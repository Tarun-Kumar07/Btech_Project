`timescale 1ns / 1ps
module convo_tb;

reg clock;
   reg reset;
    reg [24:0] in [1:0][127:0][127:0];
    reg [34:0] filter [7:0][4:0][4:0];
    reg [34:0] filter2 [31:0][4:0][4:0];
    reg [34:0] filter3 [63:0][2:0][2:0];
    reg [34:0] filter4 [127:0][2:0][2:0];
    reg [34:0] filter5 [10:0][1023:0];
    reg [34:0] bias[3:0];
    reg [34:0] bias2 [7:0];
    reg [34:0] bias3 [7:0];
    reg [34:0] bias4 [15:0];
    reg [34:0] bias5 [10:0];
    reg [7:0] pred_in [10:0];
    reg [34:0] vmem_in [3:0][63:0][63:0];
    reg [34:0] vmem_in2 [7:0][31:0][31:0];
    reg [34:0] vmem_in3 [7:0][15:0][15:0];
    reg [34:0] vmem_in4 [15:0][7:0][7:0];
    reg [34:0] vmem_in5 [10:0];
    wire [34:0] vmem_out [3:0][63:0][63:0];
    wire [34:0] vmem_out2 [7:0][31:0][31:0];
    wire [34:0] vmem_out3 [7:0][15:0][15:0];
    wire [34:0] vmem_out4 [15:0][7:0][7:0];
    reg [34:0] vmem_out5 [10:0];
    wire [7:0] pred_out[10:0];
    reg go;
    int i,j,k,t;
//    int fd;

//    reg [3:0] stride;
    wire out[3:0][63:0][63:0];
    reg [24:0]weight;
    
    int    fd, status;
  logic [15:0] mem [15:0];
  logic [34:0] reg1;
    
//layer1 l1(go,clock,reset,bias,bias2,bias3,bias4,bias5,in,filter,filter2,filter3,filter4,filter5,vmem_in,vmem_in2,vmem_in3,vmem_in4,vmem_in5, pred_in, vmem_out,vmem_out2,vmem_out3,vmem_out4,vmem_out5, pred_out);

    
    initial begin
    fd = $fopen ("values.txt", "rb");
//    $display("here");
//        bias[0]=2;
//        bias[1]=3;
//        bias[2]=1;
//        bias[3]=4;
    
//        for(int w = 0; w < 8; w++)
//        for(int i = 0; i < 5; i++)
//        for(int j = 0; j < 5; j++) begin 
//         filter[w][i][j] = 35'b00000000010100011010011111111110000;
//        end

//reg [34:0] filter [7:0][4:0][4:0];
filter[0][0][0] = 35'b11111101011001000101011010010000000;
filter[0][0][1] = 35'b00000000010100011010011111111110000;
filter[0][0][2] = 35'b11111011111001110001100101000000000;
filter[0][0][3] = 35'b00000001000111101101100010110100000;
filter[0][0][4] = 35'b00000000011001111111110010101111100;
filter[0][1][0] = 35'b11111011100101000001111111001000000;
filter[0][1][1] = 35'b11111111110000011001110001110110000;
filter[0][1][2] = 35'b00000011111010001111110010101100000;
filter[0][1][3] = 35'b11111111100001110110000111100010000;
filter[0][1][4] = 35'b11111111111100000101011110010100101;
filter[0][2][0] = 35'b11111110010110011001010000011110000;
filter[0][2][1] = 35'b00000000000101100001000000001110001;
filter[0][2][2] = 35'b11111100111010101010100100011000000;
filter[0][2][3] = 35'b00000001110001000001111001001110000;
filter[0][2][4] = 35'b11111100010101100100100110010000000;
filter[0][3][0] = 35'b00000000010101111010000011110100100;
filter[0][3][1] = 35'b00000000000000110010001110110111111;
filter[0][3][2] = 35'b00000011110011100001011011111100000;
filter[0][3][3] = 35'b00000010110110001011100000001100000;
filter[0][3][4] = 35'b11111110011000110110010000100010000;
filter[0][4][0] = 35'b11111011100010111101000001011000000;
filter[0][4][1] = 35'b11111110001011110000110110101100000;
filter[0][4][2] = 35'b00000000010110001001111000101101100;
filter[0][4][3] = 35'b00000000000011100000011010101100011;
filter[0][4][4] = 35'b00000001000111100001010100000000000;
filter[1][0][0] = 35'b00000011011111011011010101101100000;
filter[1][0][1] = 35'b11111011111011001110111001111000000;
filter[1][0][2] = 35'b11111111101010110001000111001010000;
filter[1][0][3] = 35'b00000001111100110110010000111000000;
filter[1][0][4] = 35'b11111110010111111101000001111010000;
filter[1][1][0] = 35'b00000010101000000101001110111000000;
filter[1][1][1] = 35'b11111100111100100001110101110100000;
filter[1][1][2] = 35'b00000011010011100100001000100100000;
filter[1][1][3] = 35'b11111111100000100001111011110100100;
filter[1][1][4] = 35'b00000010100101011111111000110000000;
filter[1][2][0] = 35'b11111110111011010101000111011100000;
filter[1][2][1] = 35'b11111110111011001101101010101100000;
filter[1][2][2] = 35'b00000000010111010000111001100101100;
filter[1][2][3] = 35'b00000000100011010001011011010101000;
filter[1][2][4] = 35'b00000010000100011011001110011100000;
filter[1][3][0] = 35'b11111110001011000000111000001010000;
filter[1][3][1] = 35'b00000001101111100110110010001100000;
filter[1][3][2] = 35'b11111101100101010101111100110100000;
filter[1][3][3] = 35'b11111111000111100000000011000111000;
filter[1][3][4] = 35'b11111011110001111100101101100000000;
filter[1][4][0] = 35'b11111110110010100001100111011110000;
filter[1][4][1] = 35'b11111011100000001011111010011000000;
filter[1][4][2] = 35'b11111110000101011010001100011010000;
filter[1][4][3] = 35'b11111100001000001010100010110100000;
filter[1][4][4] = 35'b11111100011111110010000011100100000;
filter[2][0][0] = 35'b00000100001010110000001100001000000;
filter[2][0][1] = 35'b00000100001001001111000001010000000;
filter[2][0][2] = 35'b00000011100110101110100011110000000;
filter[2][0][3] = 35'b11111011110011001100111110000000000;
filter[2][0][4] = 35'b11111011100001001001011001001000000;
filter[2][1][0] = 35'b00000101000110000001111110111000000;
filter[2][1][1] = 35'b11111111010001000101011100101000000;
filter[2][1][2] = 35'b11111110001001101011100001010110000;
filter[2][1][3] = 35'b11111010010110100000110010100000000;
filter[2][1][4] = 35'b11111011011101011011100100010000000;
filter[2][2][0] = 35'b00000000001001000101111101010000110;
filter[2][2][1] = 35'b11111100110110000010011100000000000;
filter[2][2][2] = 35'b11111011101000001111110011001000000;
filter[2][2][3] = 35'b11111011010110110011000011110000000;
filter[2][2][4] = 35'b11111010110010100010000100001000000;
filter[2][3][0] = 35'b00000100011100110001011111101000000;
filter[2][3][1] = 35'b00000011110001001100100101000100000;
filter[2][3][2] = 35'b11111011110000111001100000111000000;
filter[2][3][3] = 35'b00000000101101101100110100111011000;
filter[2][3][4] = 35'b11111110000011101100101110100110000;
filter[2][4][0] = 35'b11111101000000111001011100010000000;
filter[2][4][1] = 35'b00000001110101101010110110011110000;
filter[2][4][2] = 35'b11111110100011110111111010101100000;
filter[2][4][3] = 35'b11111010000001010001100110101000000;
filter[2][4][4] = 35'b00000010110000111101011110100100000;
filter[3][0][0] = 35'b00000011100100010100100011110100000;
filter[3][0][1] = 35'b00000000110101100111000111111011000;
filter[3][0][2] = 35'b11111100110100011001101010111100000;
filter[3][0][3] = 35'b11111100010111011111011010110000000;
filter[3][0][4] = 35'b11111110001010110110110110101000000;
filter[3][1][0] = 35'b00000000110111010000011000000110000;
filter[3][1][1] = 35'b11111110000011111110100010100110000;
filter[3][1][2] = 35'b00000001111010110110000100011100000;
filter[3][1][3] = 35'b11111100000111011010100100110100000;
filter[3][1][4] = 35'b00000000010010101110111110010110000;
filter[3][2][0] = 35'b11111111011100111101010010111001000;
filter[3][2][1] = 35'b00000000101001101110100011111010000;
filter[3][2][2] = 35'b11111011000001101110010111101000000;
filter[3][2][3] = 35'b11111111101011101110111101101011100;
filter[3][2][4] = 35'b11111010001101100111010000111000000;
filter[3][3][0] = 35'b11111011111100101011011000110000000;
filter[3][3][1] = 35'b00000010010100010000011111001000000;
filter[3][3][2] = 35'b11111100111010001010100011010100000;
filter[3][3][3] = 35'b11111000111011111110100101111000000;
filter[3][3][4] = 35'b11111010100000110110001111010000000;
filter[3][4][0] = 35'b00000000001101011101000000001001010;
filter[3][4][1] = 35'b00000010111101100110110111101100000;
filter[3][4][2] = 35'b11111110010011000011111011011110000;
filter[3][4][3] = 35'b11111101001000010000101000011100000;
filter[3][4][4] = 35'b11111111111101100000001101110111011;
filter[4][0][0] = 35'b11111011011111011100011100011000000;
filter[4][0][1] = 35'b00000100011101110111110000011000000;
filter[4][0][2] = 35'b11111011000000100001010010010000000;
filter[4][0][3] = 35'b11111011001011011011000101001000000;
filter[4][0][4] = 35'b11111100100011010000111111011000000;
filter[4][1][0] = 35'b11111101100010000100110100000000000;
filter[4][1][1] = 35'b00000000101110010000000001100111000;
filter[4][1][2] = 35'b11111111000110000000000100111000000;
filter[4][1][3] = 35'b00000000100011010100110001011010000;
filter[4][1][4] = 35'b11111011100001000000110000110000000;
filter[4][2][0] = 35'b11111111101101111010110010011101000;
filter[4][2][1] = 35'b00000010011111100011001010101000000;
filter[4][2][2] = 35'b00000100001001101100100110010000000;
filter[4][2][3] = 35'b00000010001101111011110111011000000;
filter[4][2][4] = 35'b11111011111101111001010010001000000;
filter[4][3][0] = 35'b11111100101101010001100010100000000;
filter[4][3][1] = 35'b11111111011111010101011111110110000;
filter[4][3][2] = 35'b11111100000101100011110010100000000;
filter[4][3][3] = 35'b11111011001000110101001110100000000;
filter[4][3][4] = 35'b11111101010011000000101110100000000;
filter[4][4][0] = 35'b00000001011110000000011010101000000;
filter[4][4][1] = 35'b00000000001110010010000100110010000;
filter[4][4][2] = 35'b00000011010110101010110111011100000;
filter[4][4][3] = 35'b11111010010111110110111110110000000;
filter[4][4][4] = 35'b11111110111101011001101000111110000;
filter[5][0][0] = 35'b11111111010001100001001001100101000;
filter[5][0][1] = 35'b00000001110011111010001000000100000;
filter[5][0][2] = 35'b11111111111110110001011011001110101;
filter[5][0][3] = 35'b11111100110100101110111010001000000;
filter[5][0][4] = 35'b11111101000001110010010101010100000;
filter[5][1][0] = 35'b00000011111010010101110111111000000;
filter[5][1][1] = 35'b11111100110000111111011001010100000;
filter[5][1][2] = 35'b00000101110101111100111101000000000;
filter[5][1][3] = 35'b00000010100011010011000010110100000;
filter[5][1][4] = 35'b11111011000011110001101001010000000;
filter[5][2][0] = 35'b11111010001001000001000100111000000;
filter[5][2][1] = 35'b00000000111010011000010000111010000;
filter[5][2][2] = 35'b00000001000000110000011110111000000;
filter[5][2][3] = 35'b11111010111010100001010110011000000;
filter[5][2][4] = 35'b11111001111010101101110111100000000;
filter[5][3][0] = 35'b11111011101010010001100000010000000;
filter[5][3][1] = 35'b11111100101100110100110110111100000;
filter[5][3][2] = 35'b00000010111000111100010010000000000;
filter[5][3][3] = 35'b11111011111000000100010001110000000;
filter[5][3][4] = 35'b11111010000001100001000111101000000;
filter[5][4][0] = 35'b00000000001101000001110001100000100;
filter[5][4][1] = 35'b11111110100011000110101001101000000;
filter[5][4][2] = 35'b00000100111111111110111111101000000;
filter[5][4][3] = 35'b11111010101101001111011100110000000;
filter[5][4][4] = 35'b11111101101011100110001100100000000;
filter[6][0][0] = 35'b11111111010110100101011110101111000;
filter[6][0][1] = 35'b00000100011111001000011010010000000;
filter[6][0][2] = 35'b00000110010111110111000011001000000;
filter[6][0][3] = 35'b00000000011101001001001100110110100;
filter[6][0][4] = 35'b00000011100111010110110000010000000;
filter[6][1][0] = 35'b00000000001000111000010000011111100;
filter[6][1][1] = 35'b00000000101111111100011100110111000;
filter[6][1][2] = 35'b00000011110010100011011001011000000;
filter[6][1][3] = 35'b00000110100000101010000000101000000;
filter[6][1][4] = 35'b11111111010010110110101111010000000;
filter[6][2][0] = 35'b11111101111001001001000001110100000;
filter[6][2][1] = 35'b00000110001000101001110110001000000;
filter[6][2][2] = 35'b00000001010101010111100001101010000;
filter[6][2][3] = 35'b11111111010111011000011010110010000;
filter[6][2][4] = 35'b00000110001101111101010000000000000;
filter[6][3][0] = 35'b00000001110010100010000110001100000;
filter[6][3][1] = 35'b00000000100000000100100011001110000;
filter[6][3][2] = 35'b00000001011001000000100001011110000;
filter[6][3][3] = 35'b00000100010000111110100111110000000;
filter[6][3][4] = 35'b00000010101101101000101100000000000;
filter[6][4][0] = 35'b11111100110101110011111100000100000;
filter[6][4][1] = 35'b00000011000110001111101111100000000;
filter[6][4][2] = 35'b00000001011000010000001001010100000;
filter[6][4][3] = 35'b00000100000111111010101101001000000;
filter[6][4][4] = 35'b00000000010110111011011011011000100;
filter[7][0][0] = 35'b00000110011100000111111101001000000;
filter[7][0][1] = 35'b00000100011111101101101011111000000;
filter[7][0][2] = 35'b11111110110111100000001001101000000;
filter[7][0][3] = 35'b11111110100000000101000111111000000;
filter[7][0][4] = 35'b11111110101011010101100001011010000;
filter[7][1][0] = 35'b00000011111010010100001110011100000;
filter[7][1][1] = 35'b00000000010110101101101110000111100;
filter[7][1][2] = 35'b00000100101111001000110100010000000;
filter[7][1][3] = 35'b00000011101111000010100110111000000;
filter[7][1][4] = 35'b00000001001110110001110000001110000;
filter[7][2][0] = 35'b00000011111010110101011000101100000;
filter[7][2][1] = 35'b11111110000001001011100010001000000;
filter[7][2][2] = 35'b00000001110100010001111101000000000;
filter[7][2][3] = 35'b11111111010010100111011001110001000;
filter[7][2][4] = 35'b00000110100001111000010110101000000;
filter[7][3][0] = 35'b00000101010011111010101110010000000;
filter[7][3][1] = 35'b11111111011110011111011101000111000;
filter[7][3][2] = 35'b11111110111110100000101110000010000;
filter[7][3][3] = 35'b00000010111000001001100000011000000;
filter[7][3][4] = 35'b00000100000000001111111101001000000;
filter[7][4][0] = 35'b00000011010100001101010100010100000;
filter[7][4][1] = 35'b11111101000110110110011100101100000;
filter[7][4][2] = 35'b00000000100011011011111000100100000;
filter[7][4][3] = 35'b00000111111010101111111000010000000;
filter[7][4][4] = 35'b00000000111001100001011000011101000;
//reg [35:0] bias [3:0];
bias[0] = 35'b11111011100110000100111101010000000;
bias[1] = 35'b00000011111000100000001000001100000;
bias[2] = 35'b00000100100000010110111110101000000;
bias[3] = 35'b00000001000010110001110101001000000;

//======================================================================


filter2[0][0][0] = 35'b00000011000011110110100111000100000;
filter2[0][0][1] = 35'b00000000110110011000110100011100000;
filter2[0][0][2] = 35'b00000010101110001101001000011000000;
filter2[0][0][3] = 35'b00000011001011111100111100101000000;
filter2[0][0][4] = 35'b11111111010100000011100000100010000;
filter2[0][1][0] = 35'b11111101110111101011111001011100000;
filter2[0][1][1] = 35'b00000000001000100010110001011111000;
filter2[0][1][2] = 35'b00000001110001111000110011110010000;
filter2[0][1][3] = 35'b00000011000011001001011000111100000;
filter2[0][1][4] = 35'b11111111110000100111001011110011110;
filter2[0][2][0] = 35'b00000010000100000000011111001000000;
filter2[0][2][1] = 35'b11111111000101001011001111110110000;
filter2[0][2][2] = 35'b00000000100011010010011110111011000;
filter2[0][2][3] = 35'b11111111000111100011100011111101000;
filter2[0][2][4] = 35'b11111101111100101000011000001000000;
filter2[0][3][0] = 35'b11111110011001001000100001111100000;
filter2[0][3][1] = 35'b00000011100010101010101111001000000;
filter2[0][3][2] = 35'b11111111010101100101011111001001000;
filter2[0][3][3] = 35'b11111101010000101110010000111100000;
filter2[0][3][4] = 35'b11111101010110110000110110100100000;
filter2[0][4][0] = 35'b00000100110100100101100111100000000;
filter2[0][4][1] = 35'b00000010001101000111000100011100000;
filter2[0][4][2] = 35'b00000010100111100010011100100100000;
filter2[0][4][3] = 35'b00000010000111101011010110110000000;
filter2[0][4][4] = 35'b00000011001001001111100010111000000;
filter2[1][0][0] = 35'b11111001111111000100011111011000000;
filter2[1][0][1] = 35'b11111001011010010011001111101000000;
filter2[1][0][2] = 35'b11111110110111000001000000110110000;
filter2[1][0][3] = 35'b11111111000011100100001011111011000;
filter2[1][0][4] = 35'b11111111100011010110101111010000000;
filter2[1][1][0] = 35'b11111000010001100010110111111000000;
filter2[1][1][1] = 35'b11111001100001100010010001100000000;
filter2[1][1][2] = 35'b11111100011010101110011111111000000;
filter2[1][1][3] = 35'b11111101100100010111001111100100000;
filter2[1][1][4] = 35'b11111010101001100010111110001000000;
filter2[1][2][0] = 35'b11111010011111101101111111101000000;
filter2[1][2][1] = 35'b11111011110010000110110100110000000;
filter2[1][2][2] = 35'b11111100011001011010111001111000000;
filter2[1][2][3] = 35'b11111010111000101101010100100000000;
filter2[1][2][4] = 35'b11111100011000010101111001110000000;
filter2[1][3][0] = 35'b11111010111100111111101001111000000;
filter2[1][3][1] = 35'b11111000001100001000011011011000000;
filter2[1][3][2] = 35'b11110111011101001011110010100000000;
filter2[1][3][3] = 35'b11111011010000110010110111101000000;
filter2[1][3][4] = 35'b11111011101111111101000000011000000;
filter2[1][4][0] = 35'b11111010111110101001011001011000000;
filter2[1][4][1] = 35'b11111010111000100010100110000000000;
filter2[1][4][2] = 35'b11110010000111000100111110110000000;
filter2[1][4][3] = 35'b11110101101011101011110010010000000;
filter2[1][4][4] = 35'b11111011011111110111010101111000000;
filter2[2][0][0] = 35'b00000000000101110111110001001000010;
filter2[2][0][1] = 35'b11111101001111110111100101000100000;
filter2[2][0][2] = 35'b11111011001111111110011011100000000;
filter2[2][0][3] = 35'b11111110011000110101110100011110000;
filter2[2][0][4] = 35'b11111111100000101001011111000100100;
filter2[2][1][0] = 35'b11111110001010100000000111011110000;
filter2[2][1][1] = 35'b11111011100011111000001111001000000;
filter2[2][1][2] = 35'b11111011011010110010000000100000000;
filter2[2][1][3] = 35'b11110111111111101100110111110000000;
filter2[2][1][4] = 35'b11111101101110111001101011011000000;
filter2[2][2][0] = 35'b11111111111001001000110000111101001;
filter2[2][2][1] = 35'b00000000001111110010111001111000110;
filter2[2][2][2] = 35'b11111001100010000100011101101000000;
filter2[2][2][3] = 35'b11111011001100101001110010011000000;
filter2[2][2][4] = 35'b11111010101101001100000011110000000;
filter2[2][3][0] = 35'b11110111010100001011111010110000000;
filter2[2][3][1] = 35'b11110111000000111011000110110000000;
filter2[2][3][2] = 35'b11110110010110111010101000100000000;
filter2[2][3][3] = 35'b11111001100101111010110001110000000;
filter2[2][3][4] = 35'b11111000011010000010111001010000000;
filter2[2][4][0] = 35'b00000000111000000011000100100110000;
filter2[2][4][1] = 35'b11111001011011000011101001110000000;
filter2[2][4][2] = 35'b11111101000000100001001011101100000;
filter2[2][4][3] = 35'b11111011010010000010110100000000000;
filter2[2][4][4] = 35'b11110111101000111010010000000000000;
filter2[3][0][0] = 35'b11111111101001010100110000111101000;
filter2[3][0][1] = 35'b00000000000100110011000001001101010;
filter2[3][0][2] = 35'b11111101001010100011001001101100000;
filter2[3][0][3] = 35'b00000000000010011111100111011000001;
filter2[3][0][4] = 35'b11111111000011011111011010111111000;
filter2[3][1][0] = 35'b11111110101000010111001110110110000;
filter2[3][1][1] = 35'b11111100100000110001110110011000000;
filter2[3][1][2] = 35'b11111111010011001011010010110010000;
filter2[3][1][3] = 35'b11111110100101110111110001000000000;
filter2[3][1][4] = 35'b11111110010101101001100101101000000;
filter2[3][2][0] = 35'b00000010001110001110101001111000000;
filter2[3][2][1] = 35'b00000011011100111110011010001100000;
filter2[3][2][2] = 35'b00000100110100101101001100011000000;
filter2[3][2][3] = 35'b00000011111101110100100011111000000;
filter2[3][2][4] = 35'b00000000100000001111000101100001000;
filter2[3][3][0] = 35'b11111111010010011000001100010001000;
filter2[3][3][1] = 35'b00000011100110000011010000001000000;
filter2[3][3][2] = 35'b00000100000010011000100000101000000;
filter2[3][3][3] = 35'b00000101000010000011010101101000000;
filter2[3][3][4] = 35'b00000101101000001101110011101000000;
filter2[3][4][0] = 35'b00000001001111001001111011011110000;
filter2[3][4][1] = 35'b11111111111110101011001111001100010;
filter2[3][4][2] = 35'b11111110001000110101100010111000000;
filter2[3][4][3] = 35'b00000100110111011001010110111000000;
filter2[3][4][4] = 35'b00000011110110001010001001010000000;
filter2[4][0][0] = 35'b11111110001100111001101001101000000;
filter2[4][0][1] = 35'b11111111000010001011011110001001000;
filter2[4][0][2] = 35'b11111111010110101010011010011100000;
filter2[4][0][3] = 35'b00000010000100010010101001010000000;
filter2[4][0][4] = 35'b00000010000001111010100000011100000;
filter2[4][1][0] = 35'b00000011011001000100100101110100000;
filter2[4][1][1] = 35'b00000000001001111101010110011100100;
filter2[4][1][2] = 35'b00000000010100110110011101101111000;
filter2[4][1][3] = 35'b00000001010100110101111111001100000;
filter2[4][1][4] = 35'b00000000111101110100110000001011000;
filter2[4][2][0] = 35'b00000001111111111111011000111010000;
filter2[4][2][1] = 35'b11111110010011011101000111100010000;
filter2[4][2][2] = 35'b00000100000111101110100100111000000;
filter2[4][2][3] = 35'b00000010011001000100100001010100000;
filter2[4][2][4] = 35'b00000010011001011000000011000100000;
filter2[4][3][0] = 35'b00000010101011011001000010011000000;
filter2[4][3][1] = 35'b00000000000110100001001001110000011;
filter2[4][3][2] = 35'b11111111001101011000011000111010000;
filter2[4][3][3] = 35'b11111111000000100011101001111101000;
filter2[4][3][4] = 35'b00000000100101011111010001111101000;
filter2[4][4][0] = 35'b11111101110000011000010000110100000;
filter2[4][4][1] = 35'b00000001011001110100011110010010000;
filter2[4][4][2] = 35'b00000010001110010111111011100100000;
filter2[4][4][3] = 35'b00000010110010010110111010110000000;
filter2[4][4][4] = 35'b00000001101011001000010011110100000;
filter2[5][0][0] = 35'b00000011000010000011011110010000000;
filter2[5][0][1] = 35'b11111110011101111101000110101000000;
filter2[5][0][2] = 35'b11111010110001111001010001010000000;
filter2[5][0][3] = 35'b00000001010010101001000011111010000;
filter2[5][0][4] = 35'b00000000111100000010110100101000000;
filter2[5][1][0] = 35'b00000010101101110010010011110100000;
filter2[5][1][1] = 35'b00000000010111100000001101100011000;
filter2[5][1][2] = 35'b11111100100001010111100001010100000;
filter2[5][1][3] = 35'b00000000000111100010111011000010000;
filter2[5][1][4] = 35'b11111011001001011111101001101000000;
filter2[5][2][0] = 35'b00000100000010110001111100100000000;
filter2[5][2][1] = 35'b11111110001101100011000110011100000;
filter2[5][2][2] = 35'b00000001011101001000110111010000000;
filter2[5][2][3] = 35'b11111111111101110010111011001111110;
filter2[5][2][4] = 35'b11111110101111000001000010001100000;
filter2[5][3][0] = 35'b11111110111010010100100100010100000;
filter2[5][3][1] = 35'b00000001101110110010110100001110000;
filter2[5][3][2] = 35'b00000100000011101110001111100000000;
filter2[5][3][3] = 35'b11111101011101101101000100100100000;
filter2[5][3][4] = 35'b11111101001010110010110101111100000;
filter2[5][4][0] = 35'b11111111111010100111100110101101001;
filter2[5][4][1] = 35'b11111110101011001000100000010100000;
filter2[5][4][2] = 35'b11111110010101001110001100111100000;
filter2[5][4][3] = 35'b00000001001001011110011101001100000;
filter2[5][4][4] = 35'b11111101110100110100001110000000000;
filter2[6][0][0] = 35'b11111111101010001011100001101101000;
filter2[6][0][1] = 35'b11111101010001101101101110000100000;
filter2[6][0][2] = 35'b11111100110101000110110010010100000;
filter2[6][0][3] = 35'b11111100000000110101010011111000000;
filter2[6][0][4] = 35'b11111100000101011001111111000100000;
filter2[6][1][0] = 35'b00000001111111100011010111000100000;
filter2[6][1][1] = 35'b11111111011011100100010010001011000;
filter2[6][1][2] = 35'b11111100101001100001000000000000000;
filter2[6][1][3] = 35'b11111101010101110001001111101000000;
filter2[6][1][4] = 35'b00000001000011001111101010100010000;
filter2[6][2][0] = 35'b11111101100100110111110110010100000;
filter2[6][2][1] = 35'b11111100011101101011100101101000000;
filter2[6][2][2] = 35'b11111110100001110100010010100010000;
filter2[6][2][3] = 35'b11111101000001101100100001010000000;
filter2[6][2][4] = 35'b00000001101100111110110010110110000;
filter2[6][3][0] = 35'b00000001111111110111111101001110000;
filter2[6][3][1] = 35'b00000001100000001001010100001000000;
filter2[6][3][2] = 35'b11111101000110100001110010011100000;
filter2[6][3][3] = 35'b00000000011001101101010111001101000;
filter2[6][3][4] = 35'b11111110100111000111110010010110000;
filter2[6][4][0] = 35'b00000100110000101110101010001000000;
filter2[6][4][1] = 35'b11111101001000000100110111001100000;
filter2[6][4][2] = 35'b00000000000010110001100010110100011;
filter2[6][4][3] = 35'b00000011100000101000110011101100000;
filter2[6][4][4] = 35'b11111011000010011101100111011000000;
filter2[7][0][0] = 35'b11111111001010001100111100010101000;
filter2[7][0][1] = 35'b00000011100110000010111000101000000;
filter2[7][0][2] = 35'b00000001011100010011001100110010000;
filter2[7][0][3] = 35'b00001000010000110001110011010000000;
filter2[7][0][4] = 35'b00001000001110011111010000110000000;
filter2[7][1][0] = 35'b11111111110110010111100101010100010;
filter2[7][1][1] = 35'b00000001101010110101010110100000000;
filter2[7][1][2] = 35'b11111111101100100110001010101100000;
filter2[7][1][3] = 35'b00000010101110000000111011010000000;
filter2[7][1][4] = 35'b00000100100010011101011000100000000;
filter2[7][2][0] = 35'b11111111000011110100101010101010000;
filter2[7][2][1] = 35'b00000000110000100000000001101100000;
filter2[7][2][2] = 35'b00000000110101001111011111011001000;
filter2[7][2][3] = 35'b00000010100001110010110010000100000;
filter2[7][2][4] = 35'b00000011101011111110010110000100000;
filter2[7][3][0] = 35'b00000001001000100011100101110000000;
filter2[7][3][1] = 35'b00000010101100100110010011111000000;
filter2[7][3][2] = 35'b00000000010111111001110111011111100;
filter2[7][3][3] = 35'b11111111010110110000111111010000000;
filter2[7][3][4] = 35'b00000000000001000101010110001001111;
filter2[7][4][0] = 35'b11111111010101110100011100011001000;
filter2[7][4][1] = 35'b11111110101010000110000100111100000;
filter2[7][4][2] = 35'b00000010111100000101100110001100000;
filter2[7][4][3] = 35'b00000001100110001000111000011110000;
filter2[7][4][4] = 35'b00000010111101100011100110110000000;
filter2[8][0][0] = 35'b11111110011011101101010100001010000;
filter2[8][0][1] = 35'b00000001010010010100010110001000000;
filter2[8][0][2] = 35'b11111111001110011010100111110101000;
filter2[8][0][3] = 35'b00000000100010000001110101111101000;
filter2[8][0][4] = 35'b11111100000101011010100101100100000;
filter2[8][1][0] = 35'b00000000100000101100001110011011000;
filter2[8][1][1] = 35'b11111101100010010000111100110000000;
filter2[8][1][2] = 35'b11111101111001110100110111101000000;
filter2[8][1][3] = 35'b11111110010001110000000011100100000;
filter2[8][1][4] = 35'b11111100011001111111011000100100000;
filter2[8][2][0] = 35'b11111101100111001101001000100100000;
filter2[8][2][1] = 35'b11111100110100110111111010011100000;
filter2[8][2][2] = 35'b11111110100000100000111110111100000;
filter2[8][2][3] = 35'b11111011010000000000000111011000000;
filter2[8][2][4] = 35'b00000001100101000100001001101010000;
filter2[8][3][0] = 35'b11111101111000011010001000110100000;
filter2[8][3][1] = 35'b11111110011100111111110001001100000;
filter2[8][3][2] = 35'b00000001001000000100101101000010000;
filter2[8][3][3] = 35'b11111101110111001101001011101000000;
filter2[8][3][4] = 35'b11111111001111110010110001011001000;
filter2[8][4][0] = 35'b11111110001000000100101101001100000;
filter2[8][4][1] = 35'b11111111001101100010100111101010000;
filter2[8][4][2] = 35'b11111011111011011100110000001000000;
filter2[8][4][3] = 35'b11111011110111011100111110110000000;
filter2[8][4][4] = 35'b11111110010100110110000001110010000;
filter2[9][0][0] = 35'b00000001100100000110110111110010000;
filter2[9][0][1] = 35'b11111101101010000011010010111100000;
filter2[9][0][2] = 35'b11111111010101101101011110100010000;
filter2[9][0][3] = 35'b11111111011110111101100100001010000;
filter2[9][0][4] = 35'b11111111111000011111010011010100100;
filter2[9][1][0] = 35'b11111110001010110000000000001110000;
filter2[9][1][1] = 35'b11111110001111110110110011111000000;
filter2[9][1][2] = 35'b00000000011001110010001111111010100;
filter2[9][1][3] = 35'b11111110011001101100001100000100000;
filter2[9][1][4] = 35'b11111100000010101100000000010100000;
filter2[9][2][0] = 35'b11111010000010101111000100110000000;
filter2[9][2][1] = 35'b11111101101110101101100010011100000;
filter2[9][2][2] = 35'b11111001111111101100111001100000000;
filter2[9][2][3] = 35'b11111100100100111111000001100100000;
filter2[9][2][4] = 35'b11111110000011000011001101110110000;
filter2[9][3][0] = 35'b11111111101101101001110011100011000;
filter2[9][3][1] = 35'b11111110010011010111000010010010000;
filter2[9][3][2] = 35'b11111010011001101111010011111000000;
filter2[9][3][3] = 35'b11111101110101100010100111110100000;
filter2[9][3][4] = 35'b00000001110110000001111001110100000;
filter2[9][4][0] = 35'b00000000110100000100110111010000000;
filter2[9][4][1] = 35'b11111111111111110000010011001001111;
filter2[9][4][2] = 35'b11111101111111010100111011010100000;
filter2[9][4][3] = 35'b11111111101011000001110001111101000;
filter2[9][4][4] = 35'b00000001110000111001110010001100000;
filter2[10][0][0] = 35'b00000000010010010101010100010000000;
filter2[10][0][1] = 35'b11111100111111110011001111000100000;
filter2[10][0][2] = 35'b11111110101000100100011110101010000;
filter2[10][0][3] = 35'b11111111001100100111110100000011000;
filter2[10][0][4] = 35'b11111111111110001111111100011101100;
filter2[10][1][0] = 35'b11111011010110101011110101000000000;
filter2[10][1][1] = 35'b11111111011001011001010010101111000;
filter2[10][1][2] = 35'b11111110111111001010001011000010000;
filter2[10][1][3] = 35'b11111011100000010111110011011000000;
filter2[10][1][4] = 35'b11111100101110010110000000011100000;
filter2[10][2][0] = 35'b00000000110000011011110011011010000;
filter2[10][2][1] = 35'b11111110000001110001001011011010000;
filter2[10][2][2] = 35'b11111001101100010110101010100000000;
filter2[10][2][3] = 35'b11111111111111110000111100010100100;
filter2[10][2][4] = 35'b11111100101011101001111111001100000;
filter2[10][3][0] = 35'b11111101011101100001100000000100000;
filter2[10][3][1] = 35'b00000000101111000001101101010011000;
filter2[10][3][2] = 35'b11111111011010100100110001010000000;
filter2[10][3][3] = 35'b11111101101101110101000011101100000;
filter2[10][3][4] = 35'b11111011011000111111111110011000000;
filter2[10][4][0] = 35'b00000000001101010110001010101111110;
filter2[10][4][1] = 35'b11111011111110111111010001110000000;
filter2[10][4][2] = 35'b00000000011001101100101111110010100;
filter2[10][4][3] = 35'b11111010110111011100101000001000000;
filter2[10][4][4] = 35'b11111100110111111111010111111000000;
filter2[11][0][0] = 35'b11111101111101101011010010110100000;
filter2[11][0][1] = 35'b00000010100001101110010111111000000;
filter2[11][0][2] = 35'b00000001011011000010100101000110000;
filter2[11][0][3] = 35'b00000010000111100100011100111100000;
filter2[11][0][4] = 35'b00000010110010001100110001001000000;
filter2[11][1][0] = 35'b00000001010101100101110001000000000;
filter2[11][1][1] = 35'b00000010000101100100000111011000000;
filter2[11][1][2] = 35'b00000110001000010010100011010000000;
filter2[11][1][3] = 35'b00000100101001000000001010011000000;
filter2[11][1][4] = 35'b00000100111111111110101110001000000;
filter2[11][2][0] = 35'b00001000110001001010100110000000000;
filter2[11][2][1] = 35'b00000110101010100101010011100000000;
filter2[11][2][2] = 35'b00000011111000011100011111110100000;
filter2[11][2][3] = 35'b00000101010101001000011101010000000;
filter2[11][2][4] = 35'b00000010000011101100000110001100000;
filter2[11][3][0] = 35'b00000101000010010110100110110000000;
filter2[11][3][1] = 35'b00000101001011111011111101000000000;
filter2[11][3][2] = 35'b00001010001000111110001100100000000;
filter2[11][3][3] = 35'b00000101001000000000100100011000000;
filter2[11][3][4] = 35'b00000100001010010100110010110000000;
filter2[11][4][0] = 35'b00000011000101110001100100011100000;
filter2[11][4][1] = 35'b00000011010001100010000011101100000;
filter2[11][4][2] = 35'b00000111100001001101010111101000000;
filter2[11][4][3] = 35'b00001001011100000100100010010000000;
filter2[11][4][4] = 35'b00000100011011100111000010000000000;
filter2[12][0][0] = 35'b11111101000000101001101111011000000;
filter2[12][0][1] = 35'b00000001000011010100001101000010000;
filter2[12][0][2] = 35'b11111100100101001010110110100000000;
filter2[12][0][3] = 35'b00000011101001000001001110111100000;
filter2[12][0][4] = 35'b00000010100010101100111100000000000;
filter2[12][1][0] = 35'b11111110100010010100100110000010000;
filter2[12][1][1] = 35'b00000001001010010101011101010000000;
filter2[12][1][2] = 35'b11111110010011000110110100100010000;
filter2[12][1][3] = 35'b00000000110111100111000101000110000;
filter2[12][1][4] = 35'b00000001000111101101010000101110000;
filter2[12][2][0] = 35'b00000000011011100010100011011111000;
filter2[12][2][1] = 35'b11111111111110111110011011001100001;
filter2[12][2][2] = 35'b00000011011001101100000111101100000;
filter2[12][2][3] = 35'b11111111110000010100100101011101000;
filter2[12][2][4] = 35'b11111101111111111001000000111000000;
filter2[12][3][0] = 35'b00000000101011101000110000101100000;
filter2[12][3][1] = 35'b11111110111000000010101110101110000;
filter2[12][3][2] = 35'b11111101101001100001101000100000000;
filter2[12][3][3] = 35'b00000000101000100011000111111001000;
filter2[12][3][4] = 35'b11111111001010001000000011010100000;
filter2[12][4][0] = 35'b11111111011110111100100001100101000;
filter2[12][4][1] = 35'b00000000000110010100010001100000100;
filter2[12][4][2] = 35'b00000011010110001001110001000100000;
filter2[12][4][3] = 35'b11111111100000110100101011010010000;
filter2[12][4][4] = 35'b00000010100001100110100100110100000;
filter2[13][0][0] = 35'b00000001001011001000111110110100000;
filter2[13][0][1] = 35'b11111101000001111101011000111000000;
filter2[13][0][2] = 35'b11111110000111001001101011101110000;
filter2[13][0][3] = 35'b11111111001010101001110010001000000;
filter2[13][0][4] = 35'b11111110110001011011010011010100000;
filter2[13][1][0] = 35'b11111101010000010111010011011000000;
filter2[13][1][1] = 35'b00000000101100111011101011110001000;
filter2[13][1][2] = 35'b11111111010110101100111100011101000;
filter2[13][1][3] = 35'b11111111010101010001111100000110000;
filter2[13][1][4] = 35'b11111110111011000001100011101010000;
filter2[13][2][0] = 35'b11111011000000010000000010010000000;
filter2[13][2][1] = 35'b00000011000010111111100111100000000;
filter2[13][2][2] = 35'b00000011011001000010001100011000000;
filter2[13][2][3] = 35'b00000001110100110100111001110000000;
filter2[13][2][4] = 35'b11111111100101100010010000111010100;
filter2[13][3][0] = 35'b11111111101111101000110110010100000;
filter2[13][3][1] = 35'b00000001001111011001010011011100000;
filter2[13][3][2] = 35'b00000010110101000001010001000000000;
filter2[13][3][3] = 35'b11111111000000001011100011110110000;
filter2[13][3][4] = 35'b11111011100110001110100000001000000;
filter2[13][4][0] = 35'b00000010111001111100111110100000000;
filter2[13][4][1] = 35'b11111111100010111111111100111110000;
filter2[13][4][2] = 35'b00000001001110110100001011110000000;
filter2[13][4][3] = 35'b00000000011110101001111100110101100;
filter2[13][4][4] = 35'b11111011001101100000011111011000000;
filter2[14][0][0] = 35'b11111111100101111110110011011010000;
filter2[14][0][1] = 35'b00000000011101010001111001111100100;
filter2[14][0][2] = 35'b11111110100000010100100100110110000;
filter2[14][0][3] = 35'b11111110001100010011011010111100000;
filter2[14][0][4] = 35'b00000001011001110000100000100110000;
filter2[14][1][0] = 35'b11111001010100001000011000101000000;
filter2[14][1][1] = 35'b00000010010001100101111110111000000;
filter2[14][1][2] = 35'b00000001100101000000011101001110000;
filter2[14][1][3] = 35'b11111110100111001001001011001110000;
filter2[14][1][4] = 35'b11111110010000010100100000011110000;
filter2[14][2][0] = 35'b11111111111100100010100011010000100;
filter2[14][2][1] = 35'b11111101110000111000001110001000000;
filter2[14][2][2] = 35'b11111100000111111110010100000000000;
filter2[14][2][3] = 35'b00000001001001000010000110011000000;
filter2[14][2][4] = 35'b00000000111101010001010110100010000;
filter2[14][3][0] = 35'b00000011111001000111111101110000000;
filter2[14][3][1] = 35'b11111110100110110001110111010110000;
filter2[14][3][2] = 35'b11111101011110000110100010001100000;
filter2[14][3][3] = 35'b00000000111000101100101001100100000;
filter2[14][3][4] = 35'b00000000001101110001100101101011110;
filter2[14][4][0] = 35'b11111100001000100010010101101000000;
filter2[14][4][1] = 35'b00000001101011010000000011011010000;
filter2[14][4][2] = 35'b00000100011110110110101101001000000;
filter2[14][4][3] = 35'b11111111000010001101101110110110000;
filter2[14][4][4] = 35'b11111110100100101111001010000100000;
filter2[15][0][0] = 35'b00000110101100101010110010100000000;
filter2[15][0][1] = 35'b11111110110010100111111100111100000;
filter2[15][0][2] = 35'b11111111100011011100010111011100000;
filter2[15][0][3] = 35'b11111101010011001010011100111000000;
filter2[15][0][4] = 35'b11111110000101101101110001111100000;
filter2[15][1][0] = 35'b00000110011011010100101000011000000;
filter2[15][1][1] = 35'b00000001000001110011001111000100000;
filter2[15][1][2] = 35'b11111111111101010000111010011000100;
filter2[15][1][3] = 35'b11111011100100001001111010011000000;
filter2[15][1][4] = 35'b11111101011111100111000010000000000;
filter2[15][2][0] = 35'b00000100100111000111001101101000000;
filter2[15][2][1] = 35'b00000101000001011111100000001000000;
filter2[15][2][2] = 35'b11111100101100111110001000001100000;
filter2[15][2][3] = 35'b11111000101110000110100011001000000;
filter2[15][2][4] = 35'b11111011110011010101101110101000000;
filter2[15][3][0] = 35'b00000001011001011011100011110000000;
filter2[15][3][1] = 35'b11111111100000011101101111111111100;
filter2[15][3][2] = 35'b11111110100000100101110000000000000;
filter2[15][3][3] = 35'b00000000000001100010100111110110100;
filter2[15][3][4] = 35'b11111111010110100111101100110001000;
filter2[15][4][0] = 35'b00000001110000100011000111010100000;
filter2[15][4][1] = 35'b00000000011000001110111001000111000;
filter2[15][4][2] = 35'b00000010001101110000010011011100000;
filter2[15][4][3] = 35'b00000000101000110111000001010001000;
filter2[15][4][4] = 35'b11111011010100011011010000101000000;
filter2[16][0][0] = 35'b11111111100011110101000011011101100;
filter2[16][0][1] = 35'b11111111001100010010100000011110000;
filter2[16][0][2] = 35'b00000010111011001111111111111100000;
filter2[16][0][3] = 35'b00000001010001001000101000111110000;
filter2[16][0][4] = 35'b11111110100000001011010000000010000;
filter2[16][1][0] = 35'b00000010000000110011000001111000000;
filter2[16][1][1] = 35'b11111100010100010111110111100100000;
filter2[16][1][2] = 35'b11111100000111101010111110110000000;
filter2[16][1][3] = 35'b11111110100001101100111010011100000;
filter2[16][1][4] = 35'b00000000100110001000000000110011000;
filter2[16][2][0] = 35'b00000010011101000110011100101100000;
filter2[16][2][1] = 35'b11111110010011100001000111101000000;
filter2[16][2][2] = 35'b11111110011111100011000111001000000;
filter2[16][2][3] = 35'b11111110000111111011011101101010000;
filter2[16][2][4] = 35'b11111111010111000110111110011111000;
filter2[16][3][0] = 35'b00000010111000110101000100101100000;
filter2[16][3][1] = 35'b00000010011100110010111101110000000;
filter2[16][3][2] = 35'b11111111110011110011111110001101110;
filter2[16][3][3] = 35'b00000001100000001101100001010010000;
filter2[16][3][4] = 35'b11111111000010010101101110001101000;
filter2[16][4][0] = 35'b00000000010111111110011101101100100;
filter2[16][4][1] = 35'b00000010001111011000110110010100000;
filter2[16][4][2] = 35'b00000011001100110011010000110000000;
filter2[16][4][3] = 35'b11111111000010111101101100000001000;
filter2[16][4][4] = 35'b11111110101000011111010010101110000;
filter2[17][0][0] = 35'b11111100010001111010001000010000000;
filter2[17][0][1] = 35'b11111111001110000111010010110001000;
filter2[17][0][2] = 35'b11111001101001111011010110100000000;
filter2[17][0][3] = 35'b11111111010010011000101001011100000;
filter2[17][0][4] = 35'b11111100110110011101111011110000000;
filter2[17][1][0] = 35'b11111011100110011011010101011000000;
filter2[17][1][1] = 35'b11111101100101000001010101010000000;
filter2[17][1][2] = 35'b11111100010010001010000001111100000;
filter2[17][1][3] = 35'b11111110001111010001110010110110000;
filter2[17][1][4] = 35'b00000100110100010000011111000000000;
filter2[17][2][0] = 35'b11111000111101001000011011001000000;
filter2[17][2][1] = 35'b11111110101010000010001100011010000;
filter2[17][2][2] = 35'b11111101010011110010011001101100000;
filter2[17][2][3] = 35'b11111101111010000111100110111100000;
filter2[17][2][4] = 35'b11111101110000101011010000001100000;
filter2[17][3][0] = 35'b11111010111001101110100101101000000;
filter2[17][3][1] = 35'b11110111010010010100111101110000000;
filter2[17][3][2] = 35'b11110111101011101111011011000000000;
filter2[17][3][3] = 35'b11111100001001001001000011110000000;
filter2[17][3][4] = 35'b00000000001100100011110001010000010;
filter2[17][4][0] = 35'b11111001011011100111011010000000000;
filter2[17][4][1] = 35'b11111010110011011111000101001000000;
filter2[17][4][2] = 35'b11111001010000111101111001111000000;
filter2[17][4][3] = 35'b11111101001100011110110000111000000;
filter2[17][4][4] = 35'b11111111110101010010001101100110100;
filter2[18][0][0] = 35'b11111101010111100111101010001000000;
filter2[18][0][1] = 35'b11111100111010111110101100010000000;
filter2[18][0][2] = 35'b11111110101101000001000100010000000;
filter2[18][0][3] = 35'b11111110110010011101110111111110000;
filter2[18][0][4] = 35'b11111111101100111110101011000110100;
filter2[18][1][0] = 35'b11111110101001010000100110111000000;
filter2[18][1][1] = 35'b11111100100111000011101111111100000;
filter2[18][1][2] = 35'b11111111101001010111110001011111000;
filter2[18][1][3] = 35'b11111111101100111111111001010110000;
filter2[18][1][4] = 35'b00000000111111100010011100000101000;
filter2[18][2][0] = 35'b11111100011000100010101110100100000;
filter2[18][2][1] = 35'b11111100001001000101110110001100000;
filter2[18][2][2] = 35'b11111010000111100011000011100000000;
filter2[18][2][3] = 35'b11111001110110101010001111001000000;
filter2[18][2][4] = 35'b11111111011000101110011011101110000;
filter2[18][3][0] = 35'b11110111101011000010011011010000000;
filter2[18][3][1] = 35'b11110111101001001110010101110000000;
filter2[18][3][2] = 35'b11110100101100110110111010100000000;
filter2[18][3][3] = 35'b11111000101111111111101111101000000;
filter2[18][3][4] = 35'b11111000110111001000010100110000000;
filter2[18][4][0] = 35'b11111001010011011011000110010000000;
filter2[18][4][1] = 35'b11111000111111011011110001111000000;
filter2[18][4][2] = 35'b11111001110111001001100100110000000;
filter2[18][4][3] = 35'b11111101010111110011010111111100000;
filter2[18][4][4] = 35'b11111111111001111101111000010111001;
filter2[19][0][0] = 35'b11111111111111000100110111000100001;
filter2[19][0][1] = 35'b00000001000101010110100110111000000;
filter2[19][0][2] = 35'b11111111001001000011011011000001000;
filter2[19][0][3] = 35'b00000000001001001101100001111110110;
filter2[19][0][4] = 35'b11111101101100100000110101010000000;
filter2[19][1][0] = 35'b00000001000010111100101100101110000;
filter2[19][1][1] = 35'b00000000111000001101001101100101000;
filter2[19][1][2] = 35'b00000000000010001111110001101011111;
filter2[19][1][3] = 35'b00000000100001011111001101001010000;
filter2[19][1][4] = 35'b11111011111010001011110001100000000;
filter2[19][2][0] = 35'b00000011011101011110011001111000000;
filter2[19][2][1] = 35'b00000100100101100011001101000000000;
filter2[19][2][2] = 35'b11111110110001101010101101111010000;
filter2[19][2][3] = 35'b11111110011100001111100011010000000;
filter2[19][2][4] = 35'b11111110010111011010001001111100000;
filter2[19][3][0] = 35'b00000100001000010111011010001000000;
filter2[19][3][1] = 35'b00000101111001111000001011110000000;
filter2[19][3][2] = 35'b00000100111110111000000110110000000;
filter2[19][3][3] = 35'b00000101100100001101001110101000000;
filter2[19][3][4] = 35'b11111110001010111010011010011000000;
filter2[19][4][0] = 35'b00000010111000000110000111111000000;
filter2[19][4][1] = 35'b00000011011110001001000111000000000;
filter2[19][4][2] = 35'b00000001111111110110001001110010000;
filter2[19][4][3] = 35'b00000001001011111001000110100110000;
filter2[19][4][4] = 35'b11111110011101011001000000101000000;
filter2[20][0][0] = 35'b11111100101111000101001100100100000;
filter2[20][0][1] = 35'b11111101010101101110101010010000000;
filter2[20][0][2] = 35'b00000010001001011001010011101000000;
filter2[20][0][3] = 35'b00000000011001100110101000110100000;
filter2[20][0][4] = 35'b00000000000100000110010101100000110;
filter2[20][1][0] = 35'b11111110111000110111101000010000000;
filter2[20][1][1] = 35'b00000001000110101100000101111110000;
filter2[20][1][2] = 35'b11111110101001010001100011101010000;
filter2[20][1][3] = 35'b00000001101001000111000000000010000;
filter2[20][1][4] = 35'b00000010001100011111010110110100000;
filter2[20][2][0] = 35'b00000000100100010001111100011111000;
filter2[20][2][1] = 35'b11111100011100000001101101111000000;
filter2[20][2][2] = 35'b11111111100010100101100011110100000;
filter2[20][2][3] = 35'b00000000000010000000001011001001001;
filter2[20][2][4] = 35'b11111110010001101101011001011100000;
filter2[20][3][0] = 35'b11111110011100010001010110001000000;
filter2[20][3][1] = 35'b11111111011010010000000110110000000;
filter2[20][3][2] = 35'b11111101111001001000101001001000000;
filter2[20][3][3] = 35'b00000001100111111001100110110010000;
filter2[20][3][4] = 35'b11111100010010101001110111011000000;
filter2[20][4][0] = 35'b11111101000011101001001011101100000;
filter2[20][4][1] = 35'b00000010010110011100111110111000000;
filter2[20][4][2] = 35'b00000010100111110101010000110100000;
filter2[20][4][3] = 35'b11111111110011010100000001011110100;
filter2[20][4][4] = 35'b11111100110111110011110010010100000;
filter2[21][0][0] = 35'b11111110001010001011000111100110000;
filter2[21][0][1] = 35'b11111101100101111100011111110000000;
filter2[21][0][2] = 35'b11111010100100010111010101000000000;
filter2[21][0][3] = 35'b11111110110101111010011111100000000;
filter2[21][0][4] = 35'b11111101110101000000000111010100000;
filter2[21][1][0] = 35'b11111101000111011010110100101100000;
filter2[21][1][1] = 35'b11111111011011111011011101011001000;
filter2[21][1][2] = 35'b11111001010000110000011100000000000;
filter2[21][1][3] = 35'b11111110000011010001110101110010000;
filter2[21][1][4] = 35'b11111011110100111111110000001000000;
filter2[21][2][0] = 35'b11111001000111011010101111010000000;
filter2[21][2][1] = 35'b11111110100110011001100101110110000;
filter2[21][2][2] = 35'b11111000100100111111101110000000000;
filter2[21][2][3] = 35'b11111001001011100000010000000000000;
filter2[21][2][4] = 35'b11111111101011000101001111011110000;
filter2[21][3][0] = 35'b11111011010110010011110011100000000;
filter2[21][3][1] = 35'b11111011011100000001000000110000000;
filter2[21][3][2] = 35'b11110111010001100111000011110000000;
filter2[21][3][3] = 35'b11111001011111100110101110010000000;
filter2[21][3][4] = 35'b11111000000010010001010001110000000;
filter2[21][4][0] = 35'b11111011011111011100100110011000000;
filter2[21][4][1] = 35'b11111010111110000011101111100000000;
filter2[21][4][2] = 35'b11111001101000001011110110000000000;
filter2[21][4][3] = 35'b11111011110111010010001000000000000;
filter2[21][4][4] = 35'b11111110010100111100001101010110000;
filter2[22][0][0] = 35'b00000000010010110110111111111111100;
filter2[22][0][1] = 35'b11111110111011011001001000101110000;
filter2[22][0][2] = 35'b11111100110001010100001011100000000;
filter2[22][0][3] = 35'b11111100101010000000011110000100000;
filter2[22][0][4] = 35'b11111011000001010101001001101000000;
filter2[22][1][0] = 35'b11111110111100110110001101111010000;
filter2[22][1][1] = 35'b11111100001001010011101001001000000;
filter2[22][1][2] = 35'b11111111110101100010101101011010010;
filter2[22][1][3] = 35'b11111001001001111101110101010000000;
filter2[22][1][4] = 35'b11111110101111000110101101110010000;
filter2[22][2][0] = 35'b11111111010001001101101001001110000;
filter2[22][2][1] = 35'b11111101101000000111011111111000000;
filter2[22][2][2] = 35'b11111001100011010110000101000000000;
filter2[22][2][3] = 35'b11111011001010000100000000111000000;
filter2[22][2][4] = 35'b11111100100000111101101001011100000;
filter2[22][3][0] = 35'b11111111101100110010011110110000000;
filter2[22][3][1] = 35'b11111101010101000011001000010000000;
filter2[22][3][2] = 35'b11111111101110110010101100110000100;
filter2[22][3][3] = 35'b11111101011010011110101110101100000;
filter2[22][3][4] = 35'b11111110000010000101001000000010000;
filter2[22][4][0] = 35'b11111110111011111001111101110000000;
filter2[22][4][1] = 35'b11111101011111100111100111011000000;
filter2[22][4][2] = 35'b11111010101110001001111001010000000;
filter2[22][4][3] = 35'b11111101000100011011111101111100000;
filter2[22][4][4] = 35'b11111010010100111011010011111000000;
filter2[23][0][0] = 35'b00000000111010010011100110010110000;
filter2[23][0][1] = 35'b11111101110111010000100111010000000;
filter2[23][0][2] = 35'b11111111010001111001001001000100000;
filter2[23][0][3] = 35'b00000000000100001001111110010110101;
filter2[23][0][4] = 35'b00000101001001001011110011110000000;
filter2[23][1][0] = 35'b00000001000111111010001100010110000;
filter2[23][1][1] = 35'b11111101110001100000111011100000000;
filter2[23][1][2] = 35'b00000000100100000111110001110110000;
filter2[23][1][3] = 35'b00000111000101010001101010111000000;
filter2[23][1][4] = 35'b00000011101000111111100100011100000;
filter2[23][2][0] = 35'b00000001110001011110011110000100000;
filter2[23][2][1] = 35'b00000010011100101111001001110000000;
filter2[23][2][2] = 35'b00000011001110101100010010000000000;
filter2[23][2][3] = 35'b00000100011111010000011000111000000;
filter2[23][2][4] = 35'b00000100011011010101101111110000000;
filter2[23][3][0] = 35'b00000000101001111010100100111011000;
filter2[23][3][1] = 35'b00000001001111101010000000101110000;
filter2[23][3][2] = 35'b00000000111011101000011110011001000;
filter2[23][3][3] = 35'b00000100010000100101011110111000000;
filter2[23][3][4] = 35'b00000011011110001010010001110000000;
filter2[23][4][0] = 35'b11111010010011100110001101110000000;
filter2[23][4][1] = 35'b11111100010000001000111010010100000;
filter2[23][4][2] = 35'b00000001001101101010100110001100000;
filter2[23][4][3] = 35'b00000001110010110000000111011100000;
filter2[23][4][4] = 35'b11111111101110101101111000001011000;
filter2[24][0][0] = 35'b00000000111111101000000101110001000;
filter2[24][0][1] = 35'b00000010010101100001100010110100000;
filter2[24][0][2] = 35'b11111110000101001100011100010110000;
filter2[24][0][3] = 35'b00000001001111110100010010100000000;
filter2[24][0][4] = 35'b11111110110001000101111111011010000;
filter2[24][1][0] = 35'b11111111101100110100100101001011100;
filter2[24][1][1] = 35'b11111100101011100100101010000100000;
filter2[24][1][2] = 35'b11111110111001011101011101011010000;
filter2[24][1][3] = 35'b00000001101101000111001011100000000;
filter2[24][1][4] = 35'b11111111010101100010001100011010000;
filter2[24][2][0] = 35'b11111101101011010101100011010100000;
filter2[24][2][1] = 35'b11111110001011101011110010111000000;
filter2[24][2][2] = 35'b11111101111101100100111001111100000;
filter2[24][2][3] = 35'b11111110001001110100100101000100000;
filter2[24][2][4] = 35'b11111011001110011011111010001000000;
filter2[24][3][0] = 35'b11111100000100111011010000100100000;
filter2[24][3][1] = 35'b00000000011100011111110110101000000;
filter2[24][3][2] = 35'b11111110000001010001010010000110000;
filter2[24][3][3] = 35'b11111101011000011010110110101100000;
filter2[24][3][4] = 35'b00000001011011011001111100111110000;
filter2[24][4][0] = 35'b11111110000001011011000010100000000;
filter2[24][4][1] = 35'b11111100001101100001010110010000000;
filter2[24][4][2] = 35'b00000000010110110001101010110100000;
filter2[24][4][3] = 35'b11111101000110000011000001011100000;
filter2[24][4][4] = 35'b11111111100110001100100101011001100;
filter2[25][0][0] = 35'b00000000001101110001100000001001110;
filter2[25][0][1] = 35'b11111010010101000011011111100000000;
filter2[25][0][2] = 35'b11111111010011100001110111100010000;
filter2[25][0][3] = 35'b11111101111110111100000100101000000;
filter2[25][0][4] = 35'b11111110101001101010111000111110000;
filter2[25][1][0] = 35'b11111011011000110110000011100000000;
filter2[25][1][1] = 35'b11111110101101000111001100000100000;
filter2[25][1][2] = 35'b00000001011101010011100100100000000;
filter2[25][1][3] = 35'b11111111110010001100111110011010110;
filter2[25][1][4] = 35'b00000010111110100011100101011000000;
filter2[25][2][0] = 35'b11111011011000101011111111010000000;
filter2[25][2][1] = 35'b11111101001101011101111110101000000;
filter2[25][2][2] = 35'b00000000101100000111101011011011000;
filter2[25][2][3] = 35'b11111100001011010010011001110000000;
filter2[25][2][4] = 35'b00000000100110000110101000111111000;
filter2[25][3][0] = 35'b11111010110011011011001100011000000;
filter2[25][3][1] = 35'b11111110111110110101101010100010000;
filter2[25][3][2] = 35'b11111111011111110101001011010001000;
filter2[25][3][3] = 35'b11111011100110011001011110100000000;
filter2[25][3][4] = 35'b11111101100011101001111110111000000;
filter2[25][4][0] = 35'b11111100011110101000111101010000000;
filter2[25][4][1] = 35'b11111100100010111001001100111100000;
filter2[25][4][2] = 35'b11110111101000001001011100010000000;
filter2[25][4][3] = 35'b11111010001101001011011001101000000;
filter2[25][4][4] = 35'b00000010011111010011100000101100000;
filter2[26][0][0] = 35'b00000101110011000000100100011000000;
filter2[26][0][1] = 35'b11111100010001100111001111010100000;
filter2[26][0][2] = 35'b00000010101101000010101001101100000;
filter2[26][0][3] = 35'b11111010111001011010101100100000000;
filter2[26][0][4] = 35'b00000011010100100011010100001000000;
filter2[26][1][0] = 35'b11111111000010001111111100101110000;
filter2[26][1][1] = 35'b00000010010000101010100101100100000;
filter2[26][1][2] = 35'b11111111100000010110010001010110100;
filter2[26][1][3] = 35'b11111110000101110010111101011010000;
filter2[26][1][4] = 35'b11111111110000100001101011110111000;
filter2[26][2][0] = 35'b11111011001100100000100101110000000;
filter2[26][2][1] = 35'b11111100001111000111111110010100000;
filter2[26][2][2] = 35'b11111100000010100000101110100100000;
filter2[26][2][3] = 35'b00000001111001101001010110010000000;
filter2[26][2][4] = 35'b11111110001011011001011101001000000;
filter2[26][3][0] = 35'b11111100110101111010001101101000000;
filter2[26][3][1] = 35'b11111110001001111001101000001010000;
filter2[26][3][2] = 35'b11111010101010110110000001101000000;
filter2[26][3][3] = 35'b11111101001101111101011100000100000;
filter2[26][3][4] = 35'b11111110001010011100001110010100000;
filter2[26][4][0] = 35'b00000000010000100101011110000011000;
filter2[26][4][1] = 35'b11111100101001110000101100010100000;
filter2[26][4][2] = 35'b11111101000000010100001100111000000;
filter2[26][4][3] = 35'b11111011100011011110100110110000000;
filter2[26][4][4] = 35'b11111101110101111101010110101100000;
filter2[27][0][0] = 35'b11111111100001000010010010101011100;
filter2[27][0][1] = 35'b11111110101100100000010110001010000;
filter2[27][0][2] = 35'b00000000010100111010101011110011100;
filter2[27][0][3] = 35'b00000010010100100001010010101000000;
filter2[27][0][4] = 35'b00000001010011111100000010100010000;
filter2[27][1][0] = 35'b00000100011010011100000111111000000;
filter2[27][1][1] = 35'b00000001000101010111010110001010000;
filter2[27][1][2] = 35'b00000101011000011011010000100000000;
filter2[27][1][3] = 35'b00000100111010001100101011101000000;
filter2[27][1][4] = 35'b00000000001101100100100011100111100;
filter2[27][2][0] = 35'b00000011111100001000101010110000000;
filter2[27][2][1] = 35'b00000010010110101111011000010000000;
filter2[27][2][2] = 35'b00000100011110110100100100100000000;
filter2[27][2][3] = 35'b00000100010001101100101101010000000;
filter2[27][2][4] = 35'b00000011110111011110000001000100000;
filter2[27][3][0] = 35'b00000011110010000011001011000100000;
filter2[27][3][1] = 35'b00000100000001010001011011010000000;
filter2[27][3][2] = 35'b00000111000101011001001001100000000;
filter2[27][3][3] = 35'b00000110010011001011101100101000000;
filter2[27][3][4] = 35'b00000000100000011101101110011110000;
filter2[27][4][0] = 35'b11111111110101000010011110000011100;
filter2[27][4][1] = 35'b00000100110010111000101101001000000;
filter2[27][4][2] = 35'b00000101111100011101010001110000000;
filter2[27][4][3] = 35'b00000011011011101101100110001000000;
filter2[27][4][4] = 35'b00000001010001101001101110110000000;
filter2[28][0][0] = 35'b11111110111100111011010100100100000;
filter2[28][0][1] = 35'b00000000101111110110100110011111000;
filter2[28][0][2] = 35'b11111101010100101110011100000100000;
filter2[28][0][3] = 35'b11111111101001000100111011000001000;
filter2[28][0][4] = 35'b00000001001001001111111110010100000;
filter2[28][1][0] = 35'b11111111010110101111010111101110000;
filter2[28][1][1] = 35'b00000001010100100001101100010000000;
filter2[28][1][2] = 35'b00000001110100001110000011001110000;
filter2[28][1][3] = 35'b00000001100000011010001110101010000;
filter2[28][1][4] = 35'b00000011000010101010110000001100000;
filter2[28][2][0] = 35'b00000000111010110011001110000101000;
filter2[28][2][1] = 35'b11111101000011101001000110100000000;
filter2[28][2][2] = 35'b11111100011010000111101000000100000;
filter2[28][2][3] = 35'b00000001111100111000011100011010000;
filter2[28][2][4] = 35'b00000000011001100100100011010000100;
filter2[28][3][0] = 35'b11111110000111111100011010001100000;
filter2[28][3][1] = 35'b00000100101001110010101111010000000;
filter2[28][3][2] = 35'b00000010111010011110111110101100000;
filter2[28][3][3] = 35'b11111101111100110100000100101100000;
filter2[28][3][4] = 35'b00000101010111100000001010100000000;
filter2[28][4][0] = 35'b11111110000111011100100100000000000;
filter2[28][4][1] = 35'b11111111111100011110110001010101011;
filter2[28][4][2] = 35'b00000011001001100101111101111100000;
filter2[28][4][3] = 35'b00000100001110110110010110010000000;
filter2[28][4][4] = 35'b00000001111010101100001101101100000;
filter2[29][0][0] = 35'b11111110001101000010101010100000000;
filter2[29][0][1] = 35'b00000000001100010010101010000100010;
filter2[29][0][2] = 35'b11111111001001110111011100101110000;
filter2[29][0][3] = 35'b00000100010000100001111110010000000;
filter2[29][0][4] = 35'b11111110111010111001110111100010000;
filter2[29][1][0] = 35'b00000010001001011011101100100000000;
filter2[29][1][1] = 35'b11111111001110110000011011111111000;
filter2[29][1][2] = 35'b00000100011110001111010011111000000;
filter2[29][1][3] = 35'b00000011111011010010000111001100000;
filter2[29][1][4] = 35'b00000001011010100101000111010000000;
filter2[29][2][0] = 35'b11111100111110011111000100110000000;
filter2[29][2][1] = 35'b11111101001000101110000111001100000;
filter2[29][2][2] = 35'b00000010111011100100010001110000000;
filter2[29][2][3] = 35'b00000011001001001011110100110100000;
filter2[29][2][4] = 35'b00000010110111100100001000110000000;
filter2[29][3][0] = 35'b00000001001111010010111111010110000;
filter2[29][3][1] = 35'b11111110110000011111011111000100000;
filter2[29][3][2] = 35'b11111111000010011101000101111101000;
filter2[29][3][3] = 35'b00000000010110111000010111111000000;
filter2[29][3][4] = 35'b00000011001010110111010111111000000;
filter2[29][4][0] = 35'b00000001110010110101100011101110000;
filter2[29][4][1] = 35'b11111111101101001001001010101100000;
filter2[29][4][2] = 35'b00000100001000101100100101010000000;
filter2[29][4][3] = 35'b00000011011001101100011110011000000;
filter2[29][4][4] = 35'b00000100010000101011101010110000000;
filter2[30][0][0] = 35'b00000011100001100010111111111000000;
filter2[30][0][1] = 35'b11111100111100011100101001111000000;
filter2[30][0][2] = 35'b00000011100011001110101000001100000;
filter2[30][0][3] = 35'b00000001010010010010100111010000000;
filter2[30][0][4] = 35'b00000011011100000000010010100100000;
filter2[30][1][0] = 35'b11111101100110101010010001101100000;
filter2[30][1][1] = 35'b00000011010100111110001111001000000;
filter2[30][1][2] = 35'b00000100110100110010101010011000000;
filter2[30][1][3] = 35'b00000111010110010000010011111000000;
filter2[30][1][4] = 35'b00000000011110010100100100011000000;
filter2[30][2][0] = 35'b11111110000110000010001010001100000;
filter2[30][2][1] = 35'b00000001110010011111100110111010000;
filter2[30][2][2] = 35'b00000010000111001111011011010000000;
filter2[30][2][3] = 35'b00000100011100010101101000111000000;
filter2[30][2][4] = 35'b00000100111001100110010101001000000;
filter2[30][3][0] = 35'b00000000110100101011010111101110000;
filter2[30][3][1] = 35'b11111111001010110100010101101011000;
filter2[30][3][2] = 35'b00000011111111010000110110101100000;
filter2[30][3][3] = 35'b11111111010100010110011001111001000;
filter2[30][3][4] = 35'b11111110101110101111010100100100000;
filter2[30][4][0] = 35'b11111110101111010100000100111110000;
filter2[30][4][1] = 35'b00000011101111110001100110111000000;
filter2[30][4][2] = 35'b00000011101111011100111110101100000;
filter2[30][4][3] = 35'b00000011010110010101101010100000000;
filter2[30][4][4] = 35'b00000000100111011010000001001101000;
filter2[31][0][0] = 35'b00000111001101010110101111001000000;
filter2[31][0][1] = 35'b11111110101001110110011001100110000;
filter2[31][0][2] = 35'b11111111111111100001100100100101100;
filter2[31][0][3] = 35'b11111011111100110001111010000000000;
filter2[31][0][4] = 35'b00000010110011010011000110001100000;
filter2[31][1][0] = 35'b00000110010110000100001000101000000;
filter2[31][1][1] = 35'b00000000110100111100101100111011000;
filter2[31][1][2] = 35'b00000000110101110101000010101100000;
filter2[31][1][3] = 35'b11111101001110110001010100000100000;
filter2[31][1][4] = 35'b11111100001011000111101001100100000;
filter2[31][2][0] = 35'b00000100001101110111101001011000000;
filter2[31][2][1] = 35'b11111101000001000001110011011000000;
filter2[31][2][2] = 35'b11111001111000001001110101000000000;
filter2[31][2][3] = 35'b11111111100011011010010010010101000;
filter2[31][2][4] = 35'b11111111111001101001110001100010011;
filter2[31][3][0] = 35'b11111111100101010100010001100000000;
filter2[31][3][1] = 35'b11111111011001111110101110001010000;
filter2[31][3][2] = 35'b11111010110100001010111110100000000;
filter2[31][3][3] = 35'b11111111101111001101110101011101000;
filter2[31][3][4] = 35'b11111101111100000000010111100100000;
filter2[31][4][0] = 35'b11111110001110111111001011010110000;
filter2[31][4][1] = 35'b11111111001111111100110101110110000;
filter2[31][4][2] = 35'b11111101100111101000110001001100000;
filter2[31][4][3] = 35'b00000011000000010011011111100000000;
filter2[31][4][4] = 35'b00000001101001010010111101010100000;

bias2[0] = 35'b11111011111011110011000101101000000;
bias2[1] = 35'b11111101101111110011110100100000000;
bias2[2] = 35'b00000010100000010110110100100000000;
bias2[3] = 35'b11111111000111101001101101011011000;
bias2[4] = 35'b11111100100001011011000001111000000;
bias2[5] = 35'b00000000001011001010001111111000000;
bias2[6] = 35'b11111110101110110011011001011000000;
bias2[7] = 35'b00000000010110110110101010000000000;
//======================================================================


filter3[0][0][0] = 35'b11111110110111010110101110110000000;
filter3[0][0][1] = 35'b00001010111110011110001110100000000;
filter3[0][0][2] = 35'b00001100001010100010011111000000000;
filter3[0][1][0] = 35'b00000011011011000000001101101000000;
filter3[0][1][1] = 35'b00001100001001100010111101110000000;
filter3[0][1][2] = 35'b00001101101100001011000111000000000;
filter3[0][2][0] = 35'b00001011110001101100010000100000000;
filter3[0][2][1] = 35'b00001110001111010110011110100000000;
filter3[0][2][2] = 35'b00000101010001011100001010001000000;
filter3[1][0][0] = 35'b11111110100110111000101000111100000;
filter3[1][0][1] = 35'b11111111000100101011101010000101000;
filter3[1][0][2] = 35'b00000011010010111100111001110000000;
filter3[1][1][0] = 35'b11111111000000000010101011001110000;
filter3[1][1][1] = 35'b11111011001010011010100010010000000;
filter3[1][1][2] = 35'b00000110110100001000111011010000000;
filter3[1][2][0] = 35'b00000000001101000010010101100001100;
filter3[1][2][1] = 35'b11111101110001011101011000001100000;
filter3[1][2][2] = 35'b00000011110110101110001001000100000;
filter3[2][0][0] = 35'b11111110011011010111011101000110000;
filter3[2][0][1] = 35'b11111111110101000010111100110001100;
filter3[2][0][2] = 35'b00000100000011101010100101010000000;
filter3[2][1][0] = 35'b11111101000101011010111010100000000;
filter3[2][1][1] = 35'b00000001011100111001110000111000000;
filter3[2][1][2] = 35'b00000100011100100011110011110000000;
filter3[2][2][0] = 35'b00000010100001100000010010011100000;
filter3[2][2][1] = 35'b00000011010000100010011001111000000;
filter3[2][2][2] = 35'b11111111010100100001101101011011000;
filter3[3][0][0] = 35'b11111100111011100111000101000100000;
filter3[3][0][1] = 35'b11110101101001100011111100010000000;
filter3[3][0][2] = 35'b11111100111100010010011010001000000;
filter3[3][1][0] = 35'b11111100010001011000011111000100000;
filter3[3][1][1] = 35'b11111010000000001011011001111000000;
filter3[3][1][2] = 35'b11111110010010001010010110001000000;
filter3[3][2][0] = 35'b11111101001110000011100100100000000;
filter3[3][2][1] = 35'b11111100110110100010001110010000000;
filter3[3][2][2] = 35'b11111001011011100001010010001000000;
filter3[4][0][0] = 35'b11111101010110110000111101010100000;
filter3[4][0][1] = 35'b00000101010001001111001110010000000;
filter3[4][0][2] = 35'b00001001111001101000111101110000000;
filter3[4][1][0] = 35'b00000100111010101101111010101000000;
filter3[4][1][1] = 35'b00001010101000100000111101000000000;
filter3[4][1][2] = 35'b00010001010000010101110100100000000;
filter3[4][2][0] = 35'b00000010011001111000101101101000000;
filter3[4][2][1] = 35'b00001011100001000111011100010000000;
filter3[4][2][2] = 35'b00001110111111010100011010000000000;
filter3[5][0][0] = 35'b11111100011011000100111101101000000;
filter3[5][0][1] = 35'b00001001000100101110110011100000000;
filter3[5][0][2] = 35'b00001011111101011101110110010000000;
filter3[5][1][0] = 35'b11111110011110010011011000111110000;
filter3[5][1][1] = 35'b00001110100100101001110100100000000;
filter3[5][1][2] = 35'b00010010001111011111011111100000000;
filter3[5][2][0] = 35'b00001001110110101000010010100000000;
filter3[5][2][1] = 35'b00010000100000010010001110000000000;
filter3[5][2][2] = 35'b00001000101001111110110000000000000;
filter3[6][0][0] = 35'b11111000110100000000101111001000000;
filter3[6][0][1] = 35'b11111110100001010000100011101000000;
filter3[6][0][2] = 35'b00000110011111011110011110100000000;
filter3[6][1][0] = 35'b11111001001110000011001111100000000;
filter3[6][1][1] = 35'b00000011001100100010110011011000000;
filter3[6][1][2] = 35'b00010000010011101011011111000000000;
filter3[6][2][0] = 35'b00000100100110111110100110100000000;
filter3[6][2][1] = 35'b00001010000001000100010000000000000;
filter3[6][2][2] = 35'b00000010110001001001011110110100000;
filter3[7][0][0] = 35'b11111111111110110001111010011101011;
filter3[7][0][1] = 35'b11111010100010010101011000001000000;
filter3[7][0][2] = 35'b00000000010111111000101001111011100;
filter3[7][1][0] = 35'b00000000101100100111001101001101000;
filter3[7][1][1] = 35'b00000001010011101110001011010010000;
filter3[7][1][2] = 35'b11111110100111011101101110000100000;
filter3[7][2][0] = 35'b00000000011000001010110100111001100;
filter3[7][2][1] = 35'b11111011100000000001011110001000000;
filter3[7][2][2] = 35'b11111111000000000001111010011010000;
filter3[8][0][0] = 35'b11111110011101101101011000111010000;
filter3[8][0][1] = 35'b00000001110111111010100111110010000;
filter3[8][0][2] = 35'b00000110101010111111111001111000000;
filter3[8][1][0] = 35'b00001010001000110001110001100000000;
filter3[8][1][1] = 35'b00001010111101010000111001010000000;
filter3[8][1][2] = 35'b00000011000011001001000111110100000;
filter3[8][2][0] = 35'b00000000000011001011000100111111110;
filter3[8][2][1] = 35'b00000011000100110100000011110000000;
filter3[8][2][2] = 35'b00000010000100101001101101111100000;
filter3[9][0][0] = 35'b00000000111101000001000001111010000;
filter3[9][0][1] = 35'b11111011110001000000110111000000000;
filter3[9][0][2] = 35'b11110110010011010110100010100000000;
filter3[9][1][0] = 35'b00000001100000011001011010101000000;
filter3[9][1][1] = 35'b00000000000111010011000110100001000;
filter3[9][1][2] = 35'b11111110100010010000100111010100000;
filter3[9][2][0] = 35'b00000010011001000100100111011100000;
filter3[9][2][1] = 35'b00000010111010000100011001001000000;
filter3[9][2][2] = 35'b00000011000011100011100011001000000;
filter3[10][0][0] = 35'b11111110001111011000001111001000000;
filter3[10][0][1] = 35'b11111110100100111100001111000110000;
filter3[10][0][2] = 35'b11111010100100100000000110101000000;
filter3[10][1][0] = 35'b11111100001010000110010010000000000;
filter3[10][1][1] = 35'b00000001010110110110100111000010000;
filter3[10][1][2] = 35'b11111111001111000011011011110111000;
filter3[10][2][0] = 35'b11111011001110101010101011100000000;
filter3[10][2][1] = 35'b11111100110100001110001001100000000;
filter3[10][2][2] = 35'b11111101110100110010110011100000000;
filter3[11][0][0] = 35'b00000001100101001101100100111100000;
filter3[11][0][1] = 35'b11111100110001010100010000101000000;
filter3[11][0][2] = 35'b00000011010111100111001101101000000;
filter3[11][1][0] = 35'b00000010100001111011011110111000000;
filter3[11][1][1] = 35'b00000001101101011101010001111010000;
filter3[11][1][2] = 35'b11111101001010111111000101111100000;
filter3[11][2][0] = 35'b11110111010101100011101111010000000;
filter3[11][2][1] = 35'b11111110111011100001010000010100000;
filter3[11][2][2] = 35'b11111110011001110010100011000000000;
filter3[12][0][0] = 35'b00000011010001111001110110011100000;
filter3[12][0][1] = 35'b11111110101011011100100011101100000;
filter3[12][0][2] = 35'b11111110100011000110011011000000000;
filter3[12][1][0] = 35'b00000001010100111000000010000010000;
filter3[12][1][1] = 35'b00000110011000100111100000111000000;
filter3[12][1][2] = 35'b00000001101101111010101100110110000;
filter3[12][2][0] = 35'b00000100011100011010100100100000000;
filter3[12][2][1] = 35'b00000011100001111001111000000000000;
filter3[12][2][2] = 35'b00000010100101000011001101110100000;
filter3[13][0][0] = 35'b11111011110110101001110001001000000;
filter3[13][0][1] = 35'b11111101100100111011010101001100000;
filter3[13][0][2] = 35'b00000010000100111010110110101000000;
filter3[13][1][0] = 35'b11111111110111010001010011110110110;
filter3[13][1][1] = 35'b00000000001101000111110001010111000;
filter3[13][1][2] = 35'b11111111100000011011010111000101100;
filter3[13][2][0] = 35'b00000101010101111101111010010000000;
filter3[13][2][1] = 35'b00000111100011010110011010110000000;
filter3[13][2][2] = 35'b00000001110101100101101110110000000;
filter3[14][0][0] = 35'b11111110011000011010111000110110000;
filter3[14][0][1] = 35'b11111111110000011001111100011011010;
filter3[14][0][2] = 35'b11111110100011111100011101110100000;
filter3[14][1][0] = 35'b11111111101111111110101001100011100;
filter3[14][1][1] = 35'b00000000000111101100011100111000101;
filter3[14][1][2] = 35'b00000010010010100111111011110100000;
filter3[14][2][0] = 35'b11111110001111111100010101011100000;
filter3[14][2][1] = 35'b00000001100010001010000001001100000;
filter3[14][2][2] = 35'b00000010110111011111011110110100000;
filter3[15][0][0] = 35'b11111001000111110100011000000000000;
filter3[15][0][1] = 35'b00000010111000010111101111000100000;
filter3[15][0][2] = 35'b00000010100110001011110101101000000;
filter3[15][1][0] = 35'b11111000100111101110100111001000000;
filter3[15][1][1] = 35'b11111111110110011001110100001010000;
filter3[15][1][2] = 35'b00000001000100101001110001010110000;
filter3[15][2][0] = 35'b11111000111110000110100101101000000;
filter3[15][2][1] = 35'b11111101011110001011100100000100000;
filter3[15][2][2] = 35'b11111101111101110010000101110100000;
filter3[16][0][0] = 35'b11110101011101001101111011010000000;
filter3[16][0][1] = 35'b11101110010001110010110011000000000;
filter3[16][0][2] = 35'b11101101011001001000100001100000000;
filter3[16][1][0] = 35'b11111011111100110000001001010000000;
filter3[16][1][1] = 35'b11110111000010100000001110110000000;
filter3[16][1][2] = 35'b11111000001110100101000011011000000;
filter3[16][2][0] = 35'b11111111100001100101010101110001100;
filter3[16][2][1] = 35'b11111001101110010010100000011000000;
filter3[16][2][2] = 35'b11111110101001111010110110110100000;
filter3[17][0][0] = 35'b11111110010010010011101100000100000;
filter3[17][0][1] = 35'b11111111100000011001111110011000000;
filter3[17][0][2] = 35'b11111110000000100010111001101110000;
filter3[17][1][0] = 35'b00000100010101111100011111101000000;
filter3[17][1][1] = 35'b11111111100110001101111000100111000;
filter3[17][1][2] = 35'b11111001011010100011010100110000000;
filter3[17][2][0] = 35'b00000000011110111110011111011101000;
filter3[17][2][1] = 35'b00000100001010000100100100101000000;
filter3[17][2][2] = 35'b11111111100111010001111010111101000;
filter3[18][0][0] = 35'b11111111101100001110010000001000100;
filter3[18][0][1] = 35'b11111101111101000001100100001000000;
filter3[18][0][2] = 35'b11111011110001010000100000111000000;
filter3[18][1][0] = 35'b00000101000100111011010010010000000;
filter3[18][1][1] = 35'b00000101011110111000100011111000000;
filter3[18][1][2] = 35'b11111110000010110000100010100010000;
filter3[18][2][0] = 35'b00001001101101100100001110100000000;
filter3[18][2][1] = 35'b00001100011011110011111011000000000;
filter3[18][2][2] = 35'b00000111101010110000101111110000000;
filter3[19][0][0] = 35'b00000000000110100010101000011110010;
filter3[19][0][1] = 35'b11111110000001010101000101001010000;
filter3[19][0][2] = 35'b11111110011010110011001010010100000;
filter3[19][1][0] = 35'b11111101010110111110010011111100000;
filter3[19][1][1] = 35'b11111111000000111100111011001011000;
filter3[19][1][2] = 35'b00000010011110011011001101001000000;
filter3[19][2][0] = 35'b00000110110111110011000010000000000;
filter3[19][2][1] = 35'b00000000011101000000111001001010000;
filter3[19][2][2] = 35'b00000000011001101001111011001011000;
filter3[20][0][0] = 35'b11111001011001001010111000010000000;
filter3[20][0][1] = 35'b11110001010111011101011110010000000;
filter3[20][0][2] = 35'b11111001000000011110000100100000000;
filter3[20][1][0] = 35'b11111001110000000111100001111000000;
filter3[20][1][1] = 35'b11110101011010001111010111110000000;
filter3[20][1][2] = 35'b11110101101011001111101101110000000;
filter3[20][2][0] = 35'b11111001111011101001011110101000000;
filter3[20][2][1] = 35'b11111110100101010001100000100010000;
filter3[20][2][2] = 35'b11111010111011101011110010000000000;
filter3[21][0][0] = 35'b11110111001110010101111000010000000;
filter3[21][0][1] = 35'b11111110001001100011101101101110000;
filter3[21][0][2] = 35'b11111000101000101010011011100000000;
filter3[21][1][0] = 35'b11111101100000010100000110101000000;
filter3[21][1][1] = 35'b11111010010010001011100000001000000;
filter3[21][1][2] = 35'b11110111011111001110000001110000000;
filter3[21][2][0] = 35'b11111110001000100111001010111000000;
filter3[21][2][1] = 35'b11111101110001001111110110111100000;
filter3[21][2][2] = 35'b11111010001111010000000011010000000;
filter3[22][0][0] = 35'b11111101011110101110010001100000000;
filter3[22][0][1] = 35'b11111100100111111001011101010100000;
filter3[22][0][2] = 35'b11111001001110000001001011100000000;
filter3[22][1][0] = 35'b00000000111010010100011010001111000;
filter3[22][1][1] = 35'b11111111001001110001011111101111000;
filter3[22][1][2] = 35'b11111011000100100010100010000000000;
filter3[22][2][0] = 35'b00000101111000101100111001001000000;
filter3[22][2][1] = 35'b00001001100011000000111000000000000;
filter3[22][2][2] = 35'b00000111110110011000100111011000000;
filter3[23][0][0] = 35'b00000000100010110011001100010100000;
filter3[23][0][1] = 35'b11111110110100000111010000001010000;
filter3[23][0][2] = 35'b11111100001011001001001111101000000;
filter3[23][1][0] = 35'b11111110111111011110001101110010000;
filter3[23][1][1] = 35'b11111110010100011001111001101000000;
filter3[23][1][2] = 35'b11111111000110000100000010100100000;
filter3[23][2][0] = 35'b11111101111010110010111011001100000;
filter3[23][2][1] = 35'b00000000111111110111111000001001000;
filter3[23][2][2] = 35'b00000001101011011011110100111100000;
filter3[24][0][0] = 35'b00000100000100001100001100100000000;
filter3[24][0][1] = 35'b00001000011100010000110110010000000;
filter3[24][0][2] = 35'b00000101011010010000000001001000000;
filter3[24][1][0] = 35'b00001011010100111010000001110000000;
filter3[24][1][1] = 35'b00001110001101001000100110010000000;
filter3[24][1][2] = 35'b00000101000110011110110101000000000;
filter3[24][2][0] = 35'b00000101100000010000111000100000000;
filter3[24][2][1] = 35'b00001110001101110010101111010000000;
filter3[24][2][2] = 35'b00000101001100100101001111001000000;
filter3[25][0][0] = 35'b11111001001011001011000100010000000;
filter3[25][0][1] = 35'b11111100101001010101010110001100000;
filter3[25][0][2] = 35'b11111011110101000100100010000000000;
filter3[25][1][0] = 35'b11111110001000100000010011100010000;
filter3[25][1][1] = 35'b11111101001010001100010011101000000;
filter3[25][1][2] = 35'b00000100001011111010000101101000000;
filter3[25][2][0] = 35'b11111111111011001000101011010011001;
filter3[25][2][1] = 35'b00000100010100100000110100101000000;
filter3[25][2][2] = 35'b00000001100011000110000111111100000;
filter3[26][0][0] = 35'b11111001001111000101001011001000000;
filter3[26][0][1] = 35'b00000000000001100011110010110011101;
filter3[26][0][2] = 35'b11111111011101000011011101100001000;
filter3[26][1][0] = 35'b11111101011000010100000001001000000;
filter3[26][1][1] = 35'b11111111011100101110110100010111000;
filter3[26][1][2] = 35'b11111111000100010100010001001101000;
filter3[26][2][0] = 35'b00000001111011110101101011110100000;
filter3[26][2][1] = 35'b00000010111010000100110110001000000;
filter3[26][2][2] = 35'b00000010010110010110000010111100000;
filter3[27][0][0] = 35'b11111101111011100100110111010000000;
filter3[27][0][1] = 35'b11111011101100100010000100001000000;
filter3[27][0][2] = 35'b11111101001100111100000000001100000;
filter3[27][1][0] = 35'b11110110000101111101010010010000000;
filter3[27][1][1] = 35'b00000001110110100110010101011100000;
filter3[27][1][2] = 35'b11111110010001101100110010000100000;
filter3[27][2][0] = 35'b11110101010011100001011111100000000;
filter3[27][2][1] = 35'b11111101011110011111100110110100000;
filter3[27][2][2] = 35'b00000000011100011100110100000111100;
filter3[28][0][0] = 35'b11111111010100000110010111001100000;
filter3[28][0][1] = 35'b11111110011000001011111010010000000;
filter3[28][0][2] = 35'b00000010111010110110000000000100000;
filter3[28][1][0] = 35'b00000010011010000011100000010000000;
filter3[28][1][1] = 35'b00001010111010000010001000100000000;
filter3[28][1][2] = 35'b00000110100010011111010010101000000;
filter3[28][2][0] = 35'b00000100011110001000000100101000000;
filter3[28][2][1] = 35'b00001011000100110001010001110000000;
filter3[28][2][2] = 35'b00001001010001110001010110110000000;
filter3[29][0][0] = 35'b11111101000001001001001110010100000;
filter3[29][0][1] = 35'b11111110111110010111111010011110000;
filter3[29][0][2] = 35'b11111111000011101011101111111011000;
filter3[29][1][0] = 35'b00000010111010100001111010011000000;
filter3[29][1][1] = 35'b00000100101010110111000000001000000;
filter3[29][1][2] = 35'b11111101010000011000000100000000000;
filter3[29][2][0] = 35'b00000100101100100001010111111000000;
filter3[29][2][1] = 35'b00000010010011101110100101000100000;
filter3[29][2][2] = 35'b00000101000011000011110111000000000;
filter3[30][0][0] = 35'b11111100110001101010110111110100000;
filter3[30][0][1] = 35'b11111110101000011100100101100000000;
filter3[30][0][2] = 35'b11111111010101010011111111001111000;
filter3[30][1][0] = 35'b11111010110011100010111101010000000;
filter3[30][1][1] = 35'b00000011000010111001111001010000000;
filter3[30][1][2] = 35'b00000010100010010001101100010100000;
filter3[30][2][0] = 35'b00000011010010101110011001000000000;
filter3[30][2][1] = 35'b00000011101111011110101100001100000;
filter3[30][2][2] = 35'b00000001010101111011011011011110000;
filter3[31][0][0] = 35'b11111011111110110001011001001000000;
filter3[31][0][1] = 35'b11111100111000101111010000100000000;
filter3[31][0][2] = 35'b11111110110101000011110110100010000;
filter3[31][1][0] = 35'b11111101100010011100001101110100000;
filter3[31][1][1] = 35'b11111111111001110000111110011101001;
filter3[31][1][2] = 35'b00000000100101000010101110110010000;
filter3[31][2][0] = 35'b11110011011110111111101101100000000;
filter3[31][2][1] = 35'b11111100010111000111111001101100000;
filter3[31][2][2] = 35'b11111110111000101011000100011110000;
filter3[32][0][0] = 35'b11111100001011110001100011110100000;
filter3[32][0][1] = 35'b11111111110111110010011000001010110;
filter3[32][0][2] = 35'b11111101011101001010101100010000000;
filter3[32][1][0] = 35'b00000001101010100001000101110100000;
filter3[32][1][1] = 35'b11111111100000010101100101001101000;
filter3[32][1][2] = 35'b11111111110111000011101100110100110;
filter3[32][2][0] = 35'b11111101111011100000110110101100000;
filter3[32][2][1] = 35'b00000000010111110010100010110111100;
filter3[32][2][2] = 35'b11111011111111100101000101001000000;
filter3[33][0][0] = 35'b11111001111111101110000011111000000;
filter3[33][0][1] = 35'b11111101110110111110110111001100000;
filter3[33][0][2] = 35'b11111000110110110100111101000000000;
filter3[33][1][0] = 35'b00000010000111000111100011000000000;
filter3[33][1][1] = 35'b11111100011101010000111100101000000;
filter3[33][1][2] = 35'b00000000000011110101110010110010001;
filter3[33][2][0] = 35'b00000001001010000111000000100000000;
filter3[33][2][1] = 35'b11111111001011011111000000010100000;
filter3[33][2][2] = 35'b11111111110010010010001001110011010;
filter3[34][0][0] = 35'b11111010101100110011111000001000000;
filter3[34][0][1] = 35'b11111100110101001011011111111000000;
filter3[34][0][2] = 35'b11111110011100000000000000010110000;
filter3[34][1][0] = 35'b11111101000110001100101001011100000;
filter3[34][1][1] = 35'b00001000001000110110010001010000000;
filter3[34][1][2] = 35'b00000100010110100011000011110000000;
filter3[34][2][0] = 35'b00000010000100110010011010110100000;
filter3[34][2][1] = 35'b00000000111010111000011100110110000;
filter3[34][2][2] = 35'b00000000101100000101111011010110000;
filter3[35][0][0] = 35'b11111110110001000100001011111010000;
filter3[35][0][1] = 35'b11111100100110111011101101010000000;
filter3[35][0][2] = 35'b11111110010010011011100010000000000;
filter3[35][1][0] = 35'b11111111000001001011110001001100000;
filter3[35][1][1] = 35'b11111011111011111111010110110000000;
filter3[35][1][2] = 35'b11111100000011111011111100011100000;
filter3[35][2][0] = 35'b00000000110010000001001001000100000;
filter3[35][2][1] = 35'b11111101000010001101000000010000000;
filter3[35][2][2] = 35'b00000011111011001001000100111100000;
filter3[36][0][0] = 35'b00000001001010001101111000111110000;
filter3[36][0][1] = 35'b00000001110010111000101110101110000;
filter3[36][0][2] = 35'b11111101010101011011011001011100000;
filter3[36][1][0] = 35'b11111011000101111010110010001000000;
filter3[36][1][1] = 35'b11111101011001101001010011101100000;
filter3[36][1][2] = 35'b11111100000101101000010111110100000;
filter3[36][2][0] = 35'b11111011101100011001011000000000000;
filter3[36][2][1] = 35'b00000001101001001110011100000100000;
filter3[36][2][2] = 35'b00000001011100001011111111011110000;
filter3[37][0][0] = 35'b00000000011100101110011001101011100;
filter3[37][0][1] = 35'b11111011011010001001110000111000000;
filter3[37][0][2] = 35'b11111100100111100110100100111000000;
filter3[37][1][0] = 35'b11111100111001011111101111000000000;
filter3[37][1][1] = 35'b00000011001011101011111001001000000;
filter3[37][1][2] = 35'b11111101110000101100111100111100000;
filter3[37][2][0] = 35'b11111101000110111010100101001100000;
filter3[37][2][1] = 35'b11111100101101000111001100011100000;
filter3[37][2][2] = 35'b11111111000011011100011011000000000;
filter3[38][0][0] = 35'b00000000100110001101110011000010000;
filter3[38][0][1] = 35'b11111100100001100100111111001000000;
filter3[38][0][2] = 35'b11111101010101010011011000101100000;
filter3[38][1][0] = 35'b00000001111111010001001100001010000;
filter3[38][1][1] = 35'b11111111110110110000100010011100100;
filter3[38][1][2] = 35'b11111111001110001110010110100111000;
filter3[38][2][0] = 35'b11110110000110011001100011110000000;
filter3[38][2][1] = 35'b11111100100010000001010111110000000;
filter3[38][2][2] = 35'b11111001100001111100111100111000000;
filter3[39][0][0] = 35'b11111000111000110001100001111000000;
filter3[39][0][1] = 35'b11111110001000000100101111010100000;
filter3[39][0][2] = 35'b11111101000110101010011111010100000;
filter3[39][1][0] = 35'b00000000001100110010011111000110100;
filter3[39][1][1] = 35'b00000001111010101001101011000100000;
filter3[39][1][2] = 35'b11111110001111011111100011110000000;
filter3[39][2][0] = 35'b11111111101001010010011111010000100;
filter3[39][2][1] = 35'b11111110011011010101100100000000000;
filter3[39][2][2] = 35'b00000110100010110011101101011000000;
filter3[40][0][0] = 35'b00001001010111101011010011100000000;
filter3[40][0][1] = 35'b11111111101101010001001010110110100;
filter3[40][0][2] = 35'b11111100101100101011110000000000000;
filter3[40][1][0] = 35'b00000110100000111000011101001000000;
filter3[40][1][1] = 35'b00000010010100000010011011110100000;
filter3[40][1][2] = 35'b11111111001100111001011111100010000;
filter3[40][2][0] = 35'b00001001001000011101101011010000000;
filter3[40][2][1] = 35'b00000100110101001000110101110000000;
filter3[40][2][2] = 35'b00000100011010010101111100110000000;
filter3[41][0][0] = 35'b11111101000011001001000110111100000;
filter3[41][0][1] = 35'b11111100111010010110100000010000000;
filter3[41][0][2] = 35'b00000000100100100100010000011001000;
filter3[41][1][0] = 35'b00000010111011111111001001011000000;
filter3[41][1][1] = 35'b00000010100111101111100011000100000;
filter3[41][1][2] = 35'b11111110110000001010011010101110000;
filter3[41][2][0] = 35'b11111110010100000011010110010110000;
filter3[41][2][1] = 35'b11111111011101010101101000001001000;
filter3[41][2][2] = 35'b11111010011111111011100110010000000;
filter3[42][0][0] = 35'b00000000000101001011111100000111010;
filter3[42][0][1] = 35'b11111011110000111000101111110000000;
filter3[42][0][2] = 35'b11111001010111101011111011011000000;
filter3[42][1][0] = 35'b11111101001010011111011001000000000;
filter3[42][1][1] = 35'b00000010010010010101000111000100000;
filter3[42][1][2] = 35'b11111111010000000001010011100111000;
filter3[42][2][0] = 35'b00000010010000100010001101001100000;
filter3[42][2][1] = 35'b11111111110000110100010101101000110;
filter3[42][2][2] = 35'b11111111001001101111100010000100000;
filter3[43][0][0] = 35'b00000000100000100100010000000110000;
filter3[43][0][1] = 35'b11111011101010000111110001110000000;
filter3[43][0][2] = 35'b00000010000100100111111011011000000;
filter3[43][1][0] = 35'b00000001001001001010111011111000000;
filter3[43][1][1] = 35'b11111110010001111111110011111000000;
filter3[43][1][2] = 35'b00000100001001011101011100111000000;
filter3[43][2][0] = 35'b00000010001000000110101101111000000;
filter3[43][2][1] = 35'b11111111100111100101010101100101100;
filter3[43][2][2] = 35'b11111101101101110111010100010100000;
filter3[44][0][0] = 35'b00000101101000010100111101010000000;
filter3[44][0][1] = 35'b00001011011010011111000000000000000;
filter3[44][0][2] = 35'b00000010000001011110111010010000000;
filter3[44][1][0] = 35'b00001001000010011111110101100000000;
filter3[44][1][1] = 35'b00000101010100011110111000101000000;
filter3[44][1][2] = 35'b11111111000110001100001001100010000;
filter3[44][2][0] = 35'b00001010000100111101011010010000000;
filter3[44][2][1] = 35'b00001011111000000100010001100000000;
filter3[44][2][2] = 35'b00000011010101101100000000011000000;
filter3[45][0][0] = 35'b00000110101010100001111011100000000;
filter3[45][0][1] = 35'b00000001010100111011000100100000000;
filter3[45][0][2] = 35'b00000011010110001111000011010000000;
filter3[45][1][0] = 35'b00000001100110000110111101010100000;
filter3[45][1][1] = 35'b11111110110010101000101100011110000;
filter3[45][1][2] = 35'b11111100110010111100100110111100000;
filter3[45][2][0] = 35'b00001000111010000101001001110000000;
filter3[45][2][1] = 35'b00000010001110111010111001101100000;
filter3[45][2][2] = 35'b11111100010101000000101101101100000;
filter3[46][0][0] = 35'b00000011100101100010000110011100000;
filter3[46][0][1] = 35'b11111101110110011001000011010000000;
filter3[46][0][2] = 35'b11111010010111101011011010011000000;
filter3[46][1][0] = 35'b00000010110101001101011101100000000;
filter3[46][1][1] = 35'b00000011001101110000111110111000000;
filter3[46][1][2] = 35'b11111100000110101111000011101000000;
filter3[46][2][0] = 35'b11111111111100101000001011000001000;
filter3[46][2][1] = 35'b00000010100100111100111110011000000;
filter3[46][2][2] = 35'b00000000111110100001010010010000000;
filter3[47][0][0] = 35'b11111010000011100000111011101000000;
filter3[47][0][1] = 35'b11111110001100001011100101111110000;
filter3[47][0][2] = 35'b11111111111110011101110011110011010;
filter3[47][1][0] = 35'b11111100111100101101001110100000000;
filter3[47][1][1] = 35'b11111110110111011001010110110010000;
filter3[47][1][2] = 35'b00000100010000001101010101000000000;
filter3[47][2][0] = 35'b11111011111110110100010101100000000;
filter3[47][2][1] = 35'b00000000010000000011001010010000000;
filter3[47][2][2] = 35'b11111111100101001101010000010110000;
filter3[48][0][0] = 35'b11111111100101000001110100110000100;
filter3[48][0][1] = 35'b11111110010000001000001011011110000;
filter3[48][0][2] = 35'b00000000000111011101100100110101111;
filter3[48][1][0] = 35'b00000001011011010101101100110010000;
filter3[48][1][1] = 35'b11111100001111101001010100100100000;
filter3[48][1][2] = 35'b11111000001001001000100000010000000;
filter3[48][2][0] = 35'b11111110110100101001101010100010000;
filter3[48][2][1] = 35'b11111000101101110000100110000000000;
filter3[48][2][2] = 35'b11110100100010010011011110100000000;
filter3[49][0][0] = 35'b00000111101110110110101010011000000;
filter3[49][0][1] = 35'b00000011011110110100010110101100000;
filter3[49][0][2] = 35'b11111110000000011100100000010000000;
filter3[49][1][0] = 35'b00000001010101101000100111010000000;
filter3[49][1][1] = 35'b00000011011100011101100101010100000;
filter3[49][1][2] = 35'b11111101100100110111011011001000000;
filter3[49][2][0] = 35'b00000010100101011100001100001100000;
filter3[49][2][1] = 35'b00000010101111101000010001011000000;
filter3[49][2][2] = 35'b11111100100011110000111010011000000;
filter3[50][0][0] = 35'b00000010101001011110010110001000000;
filter3[50][0][1] = 35'b00000100001101011010010001010000000;
filter3[50][0][2] = 35'b00000100101111111110011110101000000;
filter3[50][1][0] = 35'b11111100101001001010001001010100000;
filter3[50][1][1] = 35'b00000011000010000100000010010000000;
filter3[50][1][2] = 35'b11111110010000000000011101111000000;
filter3[50][2][0] = 35'b11111010011010110111011111110000000;
filter3[50][2][1] = 35'b11111110010101110011000010101000000;
filter3[50][2][2] = 35'b11111100110110111101011001101100000;
filter3[51][0][0] = 35'b11111111100110111011001100001111100;
filter3[51][0][1] = 35'b00000000100001110011100011000010000;
filter3[51][0][2] = 35'b00000011000011100010111111011000000;
filter3[51][1][0] = 35'b11110101011001010010011000100000000;
filter3[51][1][1] = 35'b11111110111101010000111101010000000;
filter3[51][1][2] = 35'b00000101100111001100100000000000000;
filter3[51][2][0] = 35'b00000000010001001000000001000000100;
filter3[51][2][1] = 35'b00000011010001011000010110100100000;
filter3[51][2][2] = 35'b00000000110110001000011010101001000;
filter3[52][0][0] = 35'b00000010100010011011111100001100000;
filter3[52][0][1] = 35'b00000001000111110100010100110000000;
filter3[52][0][2] = 35'b00000011101011110000010100101000000;
filter3[52][1][0] = 35'b11111100100011101101001111100100000;
filter3[52][1][1] = 35'b00000001010110001100011110100010000;
filter3[52][1][2] = 35'b00000011100100110011100110100000000;
filter3[52][2][0] = 35'b11111010001101100001111011100000000;
filter3[52][2][1] = 35'b11111010000111101111000100101000000;
filter3[52][2][2] = 35'b11111011000100100100110100001000000;
filter3[53][0][0] = 35'b00000011101010110010100011100100000;
filter3[53][0][1] = 35'b00000110001000001100000111111000000;
filter3[53][0][2] = 35'b00000001101010101010001010000110000;
filter3[53][1][0] = 35'b00000011010100101001101001101000000;
filter3[53][1][1] = 35'b00000001010110100011110001010100000;
filter3[53][1][2] = 35'b00000000001111110110111111000101100;
filter3[53][2][0] = 35'b11111011110001101011000001011000000;
filter3[53][2][1] = 35'b11111110100000001001110101010010000;
filter3[53][2][2] = 35'b11111111011110011010011010100010000;
filter3[54][0][0] = 35'b00000001101001101001000000001100000;
filter3[54][0][1] = 35'b00000110111010111110100100010000000;
filter3[54][0][2] = 35'b00000010101111010110101001111000000;
filter3[54][1][0] = 35'b11111110011001011111001110101110000;
filter3[54][1][1] = 35'b00000100000111011000011011001000000;
filter3[54][1][2] = 35'b11111101001110110001100100001000000;
filter3[54][2][0] = 35'b11111010110001101100110111100000000;
filter3[54][2][1] = 35'b00000000101100110110100001010111000;
filter3[54][2][2] = 35'b11111111100100001000000101010010000;
filter3[55][0][0] = 35'b11111001100011000000100111111000000;
filter3[55][0][1] = 35'b11111001110010111011000101100000000;
filter3[55][0][2] = 35'b00000000100100001000100001101001000;
filter3[55][1][0] = 35'b11111101110011110001001111001000000;
filter3[55][1][1] = 35'b11111110000000001111101100010100000;
filter3[55][1][2] = 35'b00000000000111111010110010110011101;
filter3[55][2][0] = 35'b11111111101000000110101111101111000;
filter3[55][2][1] = 35'b11111111010110010110100011011000000;
filter3[55][2][2] = 35'b11111111100001010010101000111010100;
filter3[56][0][0] = 35'b11111110110111101001000101110100000;
filter3[56][0][1] = 35'b00000101001100000011010101110000000;
filter3[56][0][2] = 35'b00010111000101011010001000100000000;
filter3[56][1][0] = 35'b00000000011011000100110111110111000;
filter3[56][1][1] = 35'b00001000011011100110111111110000000;
filter3[56][1][2] = 35'b00000101011110010101000001001000000;
filter3[56][2][0] = 35'b00000111001101000010011000100000000;
filter3[56][2][1] = 35'b00001001011011110010110101100000000;
filter3[56][2][2] = 35'b11111111000100111101111101111100000;
filter3[57][0][0] = 35'b11111111000111111010000110011001000;
filter3[57][0][1] = 35'b11111100001110001101011011001100000;
filter3[57][0][2] = 35'b11111011110111011111010101000000000;
filter3[57][1][0] = 35'b00000000101001000101100101000111000;
filter3[57][1][1] = 35'b00000001010000101001101001001010000;
filter3[57][1][2] = 35'b00000001100011001110111110011100000;
filter3[57][2][0] = 35'b11111010100111101101100111101000000;
filter3[57][2][1] = 35'b11111101111010111001111110101000000;
filter3[57][2][2] = 35'b00000100011001101010011110110000000;
filter3[58][0][0] = 35'b11111011000011110110100010000000000;
filter3[58][0][1] = 35'b00000011100111000011101100111000000;
filter3[58][0][2] = 35'b11111110101100011110011010011000000;
filter3[58][1][0] = 35'b11111111010100110000011011001011000;
filter3[58][1][1] = 35'b00000000010111011001110101011101100;
filter3[58][1][2] = 35'b00000011011100111000100100101100000;
filter3[58][2][0] = 35'b11111101100110110100010111110100000;
filter3[58][2][1] = 35'b11111101010100111111101111001000000;
filter3[58][2][2] = 35'b00000001011000101110010001000010000;
filter3[59][0][0] = 35'b11111101010100101011011111110000000;
filter3[59][0][1] = 35'b11110110000111010001010110110000000;
filter3[59][0][2] = 35'b11111100110111111010001011101000000;
filter3[59][1][0] = 35'b11111010011110011000110101101000000;
filter3[59][1][1] = 35'b00000000101011111011111000010110000;
filter3[59][1][2] = 35'b11111101000110010101010100100100000;
filter3[59][2][0] = 35'b11111000100101010010010110101000000;
filter3[59][2][1] = 35'b11111010001100101011110111011000000;
filter3[59][2][2] = 35'b00000000000000111100001101100011010;
filter3[60][0][0] = 35'b00000001111100101100000000000000000;
filter3[60][0][1] = 35'b11111110100110100010100110100100000;
filter3[60][0][2] = 35'b00000100000100100101011011011000000;
filter3[60][1][0] = 35'b00000010101100000010000000100000000;
filter3[60][1][1] = 35'b00000001000110000110100000110110000;
filter3[60][1][2] = 35'b00001110000111110100011001110000000;
filter3[60][2][0] = 35'b00000011001111000000100001000000000;
filter3[60][2][1] = 35'b00000011000101010011001011101000000;
filter3[60][2][2] = 35'b00001001101010001001100010110000000;
filter3[61][0][0] = 35'b00000011110000111100010001001000000;
filter3[61][0][1] = 35'b00000100100000001101100010111000000;
filter3[61][0][2] = 35'b00000110000010111000111010101000000;
filter3[61][1][0] = 35'b11111110101101011101101100111010000;
filter3[61][1][1] = 35'b00000111000111101110000110001000000;
filter3[61][1][2] = 35'b00010000011000110011010001000000000;
filter3[61][2][0] = 35'b00000011110101010000001100000100000;
filter3[61][2][1] = 35'b00000100111010010011110010000000000;
filter3[61][2][2] = 35'b00000101010111000101111010111000000;
filter3[62][0][0] = 35'b11111111010011000110010011001110000;
filter3[62][0][1] = 35'b11111111101001111100001110011110100;
filter3[62][0][2] = 35'b00000101110001111001110111101000000;
filter3[62][1][0] = 35'b11111100011001111000100010010000000;
filter3[62][1][1] = 35'b00000000111001011111011110001111000;
filter3[62][1][2] = 35'b00000011101100101011111011011000000;
filter3[62][2][0] = 35'b11111010111010110010011011111000000;
filter3[62][2][1] = 35'b11111111111101101010011110000110101;
filter3[62][2][2] = 35'b00000001010011010100001000000100000;
filter3[63][0][0] = 35'b11111111100000101010110101110110000;
filter3[63][0][1] = 35'b11111010001110010100000001001000000;
filter3[63][0][2] = 35'b11111011100010001000001110111000000;
filter3[63][1][0] = 35'b11111010000010010011110110000000000;
filter3[63][1][1] = 35'b11111111100011011100001000000100100;
filter3[63][1][2] = 35'b11111101011001110011011110111100000;
filter3[63][2][0] = 35'b11111100101110001101010011011100000;
filter3[63][2][1] = 35'b11111110100111010110100101110100000;
filter3[63][2][2] = 35'b11111111100111110010111001000011000;

bias3[0] = 35'b11111110010000010011001011100100000;
bias3[1] = 35'b11111111001100101100101110011101000;
bias3[2] = 35'b11111111000111001111110001011010000;
bias3[3] = 35'b11111101010011011100010111010100000;
bias3[4] = 35'b11111111100011100001001111000110000;
bias3[5] = 35'b11111010100101100110101001000000000;
bias3[6] = 35'b00000000100110110101110001111101000;
bias3[7] = 35'b11111101000100111110110010011100000;

//===============================================================


filter4[0][0][0] = 35'b11111110010100000100101101011100000;
filter4[0][0][1] = 35'b00000001010101100011101111101000000;
filter4[0][0][2] = 35'b11111010100001001001011110111000000;
filter4[0][1][0] = 35'b00000010000011101111100011110100000;
filter4[0][1][1] = 35'b00000011010110101100101111000100000;
filter4[0][1][2] = 35'b00000010100001001111011000100000000;
filter4[0][2][0] = 35'b11111111100110011010010100001000100;
filter4[0][2][1] = 35'b00000111100101101111111010100000000;
filter4[0][2][2] = 35'b11111111011111001101111001101101000;
filter4[1][0][0] = 35'b11111100010111101011000000110100000;
filter4[1][0][1] = 35'b11111011011110010011011001000000000;
filter4[1][0][2] = 35'b11111111011100110111000100101000000;
filter4[1][1][0] = 35'b11111000100010011100010000001000000;
filter4[1][1][1] = 35'b00000000001100011010001111010101010;
filter4[1][1][2] = 35'b00000011101000100111011001101100000;
filter4[1][2][0] = 35'b11110010110001001000010010110000000;
filter4[1][2][1] = 35'b11111101000100001100100101011100000;
filter4[1][2][2] = 35'b00000111111000111010101101100000000;
filter4[2][0][0] = 35'b11111011011101100001010101000000000;
filter4[2][0][1] = 35'b00000001000010101110110001011110000;
filter4[2][0][2] = 35'b00000010001000111111000110100000000;
filter4[2][1][0] = 35'b11111100111100011011110101011100000;
filter4[2][1][1] = 35'b11111110100001000010010010000010000;
filter4[2][1][2] = 35'b00001011110110110110001111000000000;
filter4[2][2][0] = 35'b00000001110100111100010001010110000;
filter4[2][2][1] = 35'b00000000101111011101110010100010000;
filter4[2][2][2] = 35'b00000000100010000100110011101111000;
filter4[3][0][0] = 35'b11111101110101011100001010010000000;
filter4[3][0][1] = 35'b00000001110010010110110111100010000;
filter4[3][0][2] = 35'b00000011000010100111011101000100000;
filter4[3][1][0] = 35'b11111010111001111101011000111000000;
filter4[3][1][1] = 35'b00000010100010001101110001111100000;
filter4[3][1][2] = 35'b00000111000010011011010000100000000;
filter4[3][2][0] = 35'b11111010011101000001111011111000000;
filter4[3][2][1] = 35'b00000010010010101110001010100100000;
filter4[3][2][2] = 35'b00000001000101011001110011100010000;
filter4[4][0][0] = 35'b11111101000100110011011010101000000;
filter4[4][0][1] = 35'b00000101000010010111111011010000000;
filter4[4][0][2] = 35'b11111110010011111010001011100010000;
filter4[4][1][0] = 35'b00000000011010011010110110110001000;
filter4[4][1][1] = 35'b00000100010010101010110100000000000;
filter4[4][1][2] = 35'b00000000100101011100101101011100000;
filter4[4][2][0] = 35'b00000001000100010001000110111110000;
filter4[4][2][1] = 35'b11111110001100101001010001001000000;
filter4[4][2][2] = 35'b11111101100011110000010100001100000;
filter4[5][0][0] = 35'b11111110011101100010110101001110000;
filter4[5][0][1] = 35'b11111101101000000101001110100000000;
filter4[5][0][2] = 35'b00000001100100011110010001111110000;
filter4[5][1][0] = 35'b11110111000011000011111010110000000;
filter4[5][1][1] = 35'b11111011000101111000010101100000000;
filter4[5][1][2] = 35'b00000011110001000101100011101100000;
filter4[5][2][0] = 35'b11110111100100001000101111110000000;
filter4[5][2][1] = 35'b11111100010011101110100101101100000;
filter4[5][2][2] = 35'b00000100000000010010001000110000000;
filter4[6][0][0] = 35'b00000000000010001011110001101101000;
filter4[6][0][1] = 35'b11111110010010011110100100110100000;
filter4[6][0][2] = 35'b11111100011100000010011100001100000;
filter4[6][1][0] = 35'b11111100101100100100010011010100000;
filter4[6][1][1] = 35'b00000011101110111001001010001100000;
filter4[6][1][2] = 35'b11110111111000010001000101110000000;
filter4[6][2][0] = 35'b00000100111111000110100100011000000;
filter4[6][2][1] = 35'b00001010000110100111100001000000000;
filter4[6][2][2] = 35'b00000011000011011111011111110100000;
filter4[7][0][0] = 35'b00000000001111000100000111000001100;
filter4[7][0][1] = 35'b00000010011000110111101010010100000;
filter4[7][0][2] = 35'b11111110100111111011110010101010000;
filter4[7][1][0] = 35'b11111110011010001101000000010000000;
filter4[7][1][1] = 35'b00000000100000111000111011001110000;
filter4[7][1][2] = 35'b11111110110111111110111010111100000;
filter4[7][2][0] = 35'b11111111111000100100101110101010101;
filter4[7][2][1] = 35'b00000100101111000111010100011000000;
filter4[7][2][2] = 35'b00000011111100001000110100011100000;
filter4[8][0][0] = 35'b11111101010111001101111001010000000;
filter4[8][0][1] = 35'b00000000110000101001010110010101000;
filter4[8][0][2] = 35'b11111111111001110000110101100001111;
filter4[8][1][0] = 35'b00000011101100100001101100011000000;
filter4[8][1][1] = 35'b00000100111110100111110100101000000;
filter4[8][1][2] = 35'b00001010011001010001011000100000000;
filter4[8][2][0] = 35'b00000011100000111001100010001100000;
filter4[8][2][1] = 35'b00000111001101010010010100110000000;
filter4[8][2][2] = 35'b00000111000010010000011010100000000;
filter4[9][0][0] = 35'b00000001010001111111001001010000000;
filter4[9][0][1] = 35'b11111000110011011010100010100000000;
filter4[9][0][2] = 35'b00000001001110011011000100001000000;
filter4[9][1][0] = 35'b11111111111101010010110011010001100;
filter4[9][1][1] = 35'b00000001000001010011000110010010000;
filter4[9][1][2] = 35'b00000101100110000101000011100000000;
filter4[9][2][0] = 35'b00000111001010001010001001001000000;
filter4[9][2][1] = 35'b00000011010000010010101001101100000;
filter4[9][2][2] = 35'b00000111000111111010011111111000000;
filter4[10][0][0] = 35'b11101110110010000010110111100000000;
filter4[10][0][1] = 35'b00000001000001100100001001110010000;
filter4[10][0][2] = 35'b00000000010011100101011001011111000;
filter4[10][1][0] = 35'b00000000111010010111100111110011000;
filter4[10][1][1] = 35'b00000100100010101111010010101000000;
filter4[10][1][2] = 35'b00000010101111101111011011011100000;
filter4[10][2][0] = 35'b00000101101010011001100010000000000;
filter4[10][2][1] = 35'b11111011111111010111110010100000000;
filter4[10][2][2] = 35'b11111010000110011100100010001000000;
filter4[11][0][0] = 35'b11111010100100010111110111110000000;
filter4[11][0][1] = 35'b11111100111100000101110010100000000;
filter4[11][0][2] = 35'b00000111111011000011110111000000000;
filter4[11][1][0] = 35'b11111111011010111001101101011001000;
filter4[11][1][1] = 35'b00000111011100110000100100000000000;
filter4[11][1][2] = 35'b00001000010101110000100011110000000;
filter4[11][2][0] = 35'b00000101000111100110001000000000000;
filter4[11][2][1] = 35'b00000000101011101001001000111100000;
filter4[11][2][2] = 35'b00000010010101101100100111110000000;
filter4[12][0][0] = 35'b11111111100101101110001100010011000;
filter4[12][0][1] = 35'b00000001100011011101011011100000000;
filter4[12][0][2] = 35'b00000010011110011010010000010000000;
filter4[12][1][0] = 35'b11111010110100001001001101111000000;
filter4[12][1][1] = 35'b11111100011001111001110001000100000;
filter4[12][1][2] = 35'b11111101010110100011110011001000000;
filter4[12][2][0] = 35'b11111011101110000100101100101000000;
filter4[12][2][1] = 35'b00000001111110000001000001111110000;
filter4[12][2][2] = 35'b11111100011010110001111001010000000;
filter4[13][0][0] = 35'b11111100001001011011100100010000000;
filter4[13][0][1] = 35'b11111111111000010011001111000000000;
filter4[13][0][2] = 35'b11111110100001000011001101010100000;
filter4[13][1][0] = 35'b11111100111100101110100100110100000;
filter4[13][1][1] = 35'b00000011110010010011110011100100000;
filter4[13][1][2] = 35'b00000100110110010111001010000000000;
filter4[13][2][0] = 35'b00001001011010001000000101010000000;
filter4[13][2][1] = 35'b00000011110000001011010111111000000;
filter4[13][2][2] = 35'b00001100101111100100010000010000000;
filter4[14][0][0] = 35'b00000001001000100101001110110010000;
filter4[14][0][1] = 35'b11111100110111101101101001111000000;
filter4[14][0][2] = 35'b00000000100110100010001001011111000;
filter4[14][1][0] = 35'b11110110011100000001001011010000000;
filter4[14][1][1] = 35'b11111101100101100000101111110000000;
filter4[14][1][2] = 35'b00000011101011000110110001100000000;
filter4[14][2][0] = 35'b11111100010011010101011101100100000;
filter4[14][2][1] = 35'b00000000100110111001100000000010000;
filter4[14][2][2] = 35'b00000101010011010100110011001000000;
filter4[15][0][0] = 35'b00000001000100111110100111000100000;
filter4[15][0][1] = 35'b00000000010011010111000110110000100;
filter4[15][0][2] = 35'b00000000111010110110110100101011000;
filter4[15][1][0] = 35'b00000010100000000110101111011000000;
filter4[15][1][1] = 35'b11111111100110110110111001000101000;
filter4[15][1][2] = 35'b00000010011111010100010100100100000;
filter4[15][2][0] = 35'b11111111101010010011011100010000000;
filter4[15][2][1] = 35'b00000111111000101011111011000000000;
filter4[15][2][2] = 35'b11111101110011100000110101010000000;
filter4[16][0][0] = 35'b11111100011101011101000101111100000;
filter4[16][0][1] = 35'b11110110111011111100100001010000000;
filter4[16][0][2] = 35'b11111001011110000101001011001000000;
filter4[16][1][0] = 35'b00000000101010101111010111101111000;
filter4[16][1][1] = 35'b11111111000110111011100110100111000;
filter4[16][1][2] = 35'b00000000101111001101010001100110000;
filter4[16][2][0] = 35'b00000000110010101000011111110100000;
filter4[16][2][1] = 35'b00001000110011111000001000000000000;
filter4[16][2][2] = 35'b00000010110100110000011111101000000;
filter4[17][0][0] = 35'b00000001011001100011000000100100000;
filter4[17][0][1] = 35'b11110111011100000001011011010000000;
filter4[17][0][2] = 35'b00000000101000001111110111100001000;
filter4[17][1][0] = 35'b00000001100000011110011110001000000;
filter4[17][1][1] = 35'b00000100110110001010111010100000000;
filter4[17][1][2] = 35'b11111111101111110100101101001010000;
filter4[17][2][0] = 35'b00001010101010100100101111110000000;
filter4[17][2][1] = 35'b00000010111111000010110100101000000;
filter4[17][2][2] = 35'b00000000100111111110101010000111000;
filter4[18][0][0] = 35'b11111101110000110001100000111000000;
filter4[18][0][1] = 35'b11111100001011000001110000110000000;
filter4[18][0][2] = 35'b11111110011001001110001001001010000;
filter4[18][1][0] = 35'b00000000001100110011110011000010010;
filter4[18][1][1] = 35'b00000010100111001001111111011100000;
filter4[18][1][2] = 35'b00000000000010001001010100101000000;
filter4[18][2][0] = 35'b11111111110111001111101011101100000;
filter4[18][2][1] = 35'b00000000011010101111111101111011100;
filter4[18][2][2] = 35'b11111110011110011000000101010110000;
filter4[19][0][0] = 35'b11111000010111001100110000110000000;
filter4[19][0][1] = 35'b11110111100101110111010111100000000;
filter4[19][0][2] = 35'b11110110111100001000010111010000000;
filter4[19][1][0] = 35'b11111110001010001000000011101010000;
filter4[19][1][1] = 35'b11111110011111001000101111100110000;
filter4[19][1][2] = 35'b00000101001101011101001111100000000;
filter4[19][2][0] = 35'b00000110111111000111101001000000000;
filter4[19][2][1] = 35'b00000101010010101111000001011000000;
filter4[19][2][2] = 35'b11111110011100000101111010011100000;
filter4[20][0][0] = 35'b00000101101000101101101111110000000;
filter4[20][0][1] = 35'b11111011100011110001001011101000000;
filter4[20][0][2] = 35'b00000011010001101110111000111000000;
filter4[20][1][0] = 35'b11111110100000001000110100100100000;
filter4[20][1][1] = 35'b11111101101001000101010101101100000;
filter4[20][1][2] = 35'b11111011101101110100110010010000000;
filter4[20][2][0] = 35'b00000010001011010110001100110000000;
filter4[20][2][1] = 35'b11111110101111001000111100111110000;
filter4[20][2][2] = 35'b00000000010000001100100111011010100;
filter4[21][0][0] = 35'b00000001000010001100111000001110000;
filter4[21][0][1] = 35'b11111000111001011000101101011000000;
filter4[21][0][2] = 35'b00000010011010111011000101100000000;
filter4[21][1][0] = 35'b00000000000001110111000101110111010;
filter4[21][1][1] = 35'b00000011000100100111100110111100000;
filter4[21][1][2] = 35'b11111010101101011000111111111000000;
filter4[21][2][0] = 35'b00000011101111111011100100000000000;
filter4[21][2][1] = 35'b00000110100001101101110110011000000;
filter4[21][2][2] = 35'b11111101110011111001001011110000000;
filter4[22][0][0] = 35'b00000001111001111111000100101000000;
filter4[22][0][1] = 35'b00000000100111010001101001110001000;
filter4[22][0][2] = 35'b11111010111011111010111000001000000;
filter4[22][1][0] = 35'b11111101010001101001111011001000000;
filter4[22][1][1] = 35'b11110101011010101000011010010000000;
filter4[22][1][2] = 35'b11111000101010110001001110101000000;
filter4[22][2][0] = 35'b00000010100000001101111110010000000;
filter4[22][2][1] = 35'b11111100111011010011111001001100000;
filter4[22][2][2] = 35'b00000100101011011101100010100000000;
filter4[23][0][0] = 35'b11111010011001010110100110010000000;
filter4[23][0][1] = 35'b11111100010000001010010001101100000;
filter4[23][0][2] = 35'b11111010000001100001100111011000000;
filter4[23][1][0] = 35'b11111100000011101011100111101100000;
filter4[23][1][1] = 35'b11111100101101001010011100001100000;
filter4[23][1][2] = 35'b11111111101111110000101010011010000;
filter4[23][2][0] = 35'b00000010111111010111000101101000000;
filter4[23][2][1] = 35'b00001010001111100101100000100000000;
filter4[23][2][2] = 35'b11111111111101111010011111111111011;
filter4[24][0][0] = 35'b11111111011010000100101111010111000;
filter4[24][0][1] = 35'b00000001010101011100100011010100000;
filter4[24][0][2] = 35'b00000000011110111000000010100001000;
filter4[24][1][0] = 35'b00001001000101000111111101000000000;
filter4[24][1][1] = 35'b00000011001001010100010101111000000;
filter4[24][1][2] = 35'b11111101101010000011011011110000000;
filter4[24][2][0] = 35'b00000110000011111010111011111000000;
filter4[24][2][1] = 35'b00000010011101110010111100111100000;
filter4[24][2][2] = 35'b11111110011101111110111001011110000;
filter4[25][0][0] = 35'b00000101011001110000111010101000000;
filter4[25][0][1] = 35'b11111011011001011011011111101000000;
filter4[25][0][2] = 35'b11111111011011111111101010011110000;
filter4[25][1][0] = 35'b00000111001010111100000110011000000;
filter4[25][1][1] = 35'b00001010010110100010011000000000000;
filter4[25][1][2] = 35'b00000100010010000100011010010000000;
filter4[25][2][0] = 35'b11111011001110000100000010100000000;
filter4[25][2][1] = 35'b00000101000000000000101011001000000;
filter4[25][2][2] = 35'b11111100101110111110001100011000000;
filter4[26][0][0] = 35'b11111110001110101101001100001010000;
filter4[26][0][1] = 35'b00000110010111000000101011111000000;
filter4[26][0][2] = 35'b11110111011111101110100001000000000;
filter4[26][1][0] = 35'b11111100110111001110100101011100000;
filter4[26][1][1] = 35'b11111111110100101000111101111110100;
filter4[26][1][2] = 35'b11110110001010100111100000110000000;
filter4[26][2][0] = 35'b11111101111010111101100110011100000;
filter4[26][2][1] = 35'b11111101001000011110001100001100000;
filter4[26][2][2] = 35'b00000011011110011101011110010100000;
filter4[27][0][0] = 35'b00001001100100001001000111100000000;
filter4[27][0][1] = 35'b00000010001000101101011110111000000;
filter4[27][0][2] = 35'b11111111001111111101000100000101000;
filter4[27][1][0] = 35'b00001000001010101010101100100000000;
filter4[27][1][1] = 35'b00001001110100100001100110010000000;
filter4[27][1][2] = 35'b00000011110000001101001001011000000;
filter4[27][2][0] = 35'b11111011100000110011011001001000000;
filter4[27][2][1] = 35'b00000001110010111001011111011100000;
filter4[27][2][2] = 35'b11111100101110101100010110111100000;
filter4[28][0][0] = 35'b00000001100101000011110110010110000;
filter4[28][0][1] = 35'b11111011001100011000011101100000000;
filter4[28][0][2] = 35'b11111111000100101000100101101011000;
filter4[28][1][0] = 35'b00000001010100010111100110001100000;
filter4[28][1][1] = 35'b00000001101010101110110000010010000;
filter4[28][1][2] = 35'b00000111111000111011111101010000000;
filter4[28][2][0] = 35'b00000011101011010111011110010100000;
filter4[28][2][1] = 35'b00000001011011011100011110010110000;
filter4[28][2][2] = 35'b11111010010101101101011100000000000;
filter4[29][0][0] = 35'b00000101110111000000111000011000000;
filter4[29][0][1] = 35'b00000001010010101011101101011110000;
filter4[29][0][2] = 35'b11111100111110100001111011111000000;
filter4[29][1][0] = 35'b00000010101011001011110000100000000;
filter4[29][1][1] = 35'b00001101000101111010100010110000000;
filter4[29][1][2] = 35'b00000101101000001001001110011000000;
filter4[29][2][0] = 35'b11111010001111111111011111101000000;
filter4[29][2][1] = 35'b00000010100000010001010101111100000;
filter4[29][2][2] = 35'b11111100100101011111000011111000000;
filter4[30][0][0] = 35'b11111010101101011110010110111000000;
filter4[30][0][1] = 35'b11111000110000101011010111101000000;
filter4[30][0][2] = 35'b00000001001000110111001110011110000;
filter4[30][1][0] = 35'b00000001110011101001100101011010000;
filter4[30][1][1] = 35'b11111111011111000000110010010010000;
filter4[30][1][2] = 35'b11110110001111100010011111100000000;
filter4[30][2][0] = 35'b00000010001110000000100010100100000;
filter4[30][2][1] = 35'b11111111011010010111110100011110000;
filter4[30][2][2] = 35'b00000010111011110110000100111000000;
filter4[31][0][0] = 35'b11111101100010110100011110101100000;
filter4[31][0][1] = 35'b00000001010000111111101010000110000;
filter4[31][0][2] = 35'b00001000110000000100100000010000000;
filter4[31][1][0] = 35'b00001000010010000000000011110000000;
filter4[31][1][1] = 35'b00000000000011110011100111011010111;
filter4[31][1][2] = 35'b11111100010010100100101010111100000;
filter4[31][2][0] = 35'b00000100001110111011011110111000000;
filter4[31][2][1] = 35'b00000000101100110011110111010100000;
filter4[31][2][2] = 35'b00000000010011111010111010011000000;
filter4[32][0][0] = 35'b00000001101110101101001010110100000;
filter4[32][0][1] = 35'b11111110110001110111111100110000000;
filter4[32][0][2] = 35'b11111101001000010001100001001100000;
filter4[32][1][0] = 35'b00000000111000100010110011010111000;
filter4[32][1][1] = 35'b00000100111100110010010010101000000;
filter4[32][1][2] = 35'b00000000001101110110000011010101000;
filter4[32][2][0] = 35'b11111100111000110000001110000100000;
filter4[32][2][1] = 35'b00000000100001110111111100011010000;
filter4[32][2][2] = 35'b11111111011100111100111110101111000;
filter4[33][0][0] = 35'b11111110100010010010100110101110000;
filter4[33][0][1] = 35'b00000000110001010110110001111000000;
filter4[33][0][2] = 35'b11111110000100110011111011001110000;
filter4[33][1][0] = 35'b00000010001111110001100100011100000;
filter4[33][1][1] = 35'b00000010010001000101000011101000000;
filter4[33][1][2] = 35'b00001001101011011001010111000000000;
filter4[33][2][0] = 35'b00001010010011110011101100110000000;
filter4[33][2][1] = 35'b00000000101010010000010111011111000;
filter4[33][2][2] = 35'b00000001111010100001101110000000000;
filter4[34][0][0] = 35'b11110110001000101001110110100000000;
filter4[34][0][1] = 35'b11111011010001000111110111100000000;
filter4[34][0][2] = 35'b11111101101110000110100001010000000;
filter4[34][1][0] = 35'b11111100100100000101000111111000000;
filter4[34][1][1] = 35'b11111111110110100011101110010000010;
filter4[34][1][2] = 35'b11111110001010010111010110010010000;
filter4[34][2][0] = 35'b11110111011011100001110011110000000;
filter4[34][2][1] = 35'b11110101010010100100001000100000000;
filter4[34][2][2] = 35'b11111001111111110101100111001000000;
filter4[35][0][0] = 35'b00000000011100100001011101011011100;
filter4[35][0][1] = 35'b00000110000100100111000011000000000;
filter4[35][0][2] = 35'b11111111011010110010001000111110000;
filter4[35][1][0] = 35'b00000001101000110010010111011110000;
filter4[35][1][1] = 35'b00000010000110010111110100100000000;
filter4[35][1][2] = 35'b00000101010110110000110101010000000;
filter4[35][2][0] = 35'b00000100101100100100000011000000000;
filter4[35][2][1] = 35'b00000001111110110001010001110100000;
filter4[35][2][2] = 35'b00000100000000001101001000110000000;
filter4[36][0][0] = 35'b11111000111111010010100010100000000;
filter4[36][0][1] = 35'b11111110110011111011010001111110000;
filter4[36][0][2] = 35'b00000010111101110100110110100000000;
filter4[36][1][0] = 35'b00000101001110001100011110101000000;
filter4[36][1][1] = 35'b11111100000101100001010111000100000;
filter4[36][1][2] = 35'b11111000101001011010001000101000000;
filter4[36][2][0] = 35'b11111101001111011111001111110000000;
filter4[36][2][1] = 35'b11111111101000010110000011011101100;
filter4[36][2][2] = 35'b11111110011010011011100100011110000;
filter4[37][0][0] = 35'b00000110111010010010011100000000000;
filter4[37][0][1] = 35'b00000010111111110111111011010000000;
filter4[37][0][2] = 35'b00000100011100000111100010010000000;
filter4[37][1][0] = 35'b11111011100001010110110011000000000;
filter4[37][1][1] = 35'b00000000001100000000110011001100110;
filter4[37][1][2] = 35'b00000011110111101010111011100100000;
filter4[37][2][0] = 35'b00000111110001101001010001000000000;
filter4[37][2][1] = 35'b00000000011111001000101111000100100;
filter4[37][2][2] = 35'b11111110001101010011000110010000000;
filter4[38][0][0] = 35'b00000010000111100011101101100100000;
filter4[38][0][1] = 35'b00000011101101000001000100111100000;
filter4[38][0][2] = 35'b11110111100101010101101101010000000;
filter4[38][1][0] = 35'b11111010001011110011010101111000000;
filter4[38][1][1] = 35'b00000001110110011101111010010100000;
filter4[38][1][2] = 35'b11111100001110110111100111000000000;
filter4[38][2][0] = 35'b11110100000111001000111111010000000;
filter4[38][2][1] = 35'b11111110011001100110111110101000000;
filter4[38][2][2] = 35'b00000100111111100110100000101000000;
filter4[39][0][0] = 35'b00000110010111000000010000110000000;
filter4[39][0][1] = 35'b11111101100101100110100011111100000;
filter4[39][0][2] = 35'b11111001000010100110001001001000000;
filter4[39][1][0] = 35'b11111100110100110101011000101000000;
filter4[39][1][1] = 35'b00000100000110011111110111010000000;
filter4[39][1][2] = 35'b00000011000101001110001100111000000;
filter4[39][2][0] = 35'b11111110001010100010000010100000000;
filter4[39][2][1] = 35'b11111111000111000101100101111010000;
filter4[39][2][2] = 35'b00000100011110010001000011100000000;
filter4[40][0][0] = 35'b11111111110111110111100101010011100;
filter4[40][0][1] = 35'b11111110000010110110010110010110000;
filter4[40][0][2] = 35'b11111111101110101001011101001101100;
filter4[40][1][0] = 35'b11111111111101001110000001001100011;
filter4[40][1][1] = 35'b00000101010101101000010000001000000;
filter4[40][1][2] = 35'b11111101100110010011011100100100000;
filter4[40][2][0] = 35'b00000001101010110101111010010000000;
filter4[40][2][1] = 35'b00001110110111011010000011010000000;
filter4[40][2][2] = 35'b00000101100001000000011111010000000;
filter4[41][0][0] = 35'b11111111110010101101010110011011110;
filter4[41][0][1] = 35'b11111101010000011100101111011100000;
filter4[41][0][2] = 35'b11111100011001000100100010010000000;
filter4[41][1][0] = 35'b00000111000011110100111011010000000;
filter4[41][1][1] = 35'b00000111010011000111010110110000000;
filter4[41][1][2] = 35'b11111111110011110000111011101111010;
filter4[41][2][0] = 35'b11111011011100010100110001011000000;
filter4[41][2][1] = 35'b00000110110100111010110011000000000;
filter4[41][2][2] = 35'b11111011101001010111001001111000000;
filter4[42][0][0] = 35'b11111100001110111100000101100000000;
filter4[42][0][1] = 35'b00000110111100001000110000100000000;
filter4[42][0][2] = 35'b11111110100110011100011001110100000;
filter4[42][1][0] = 35'b11111000010100011110000011011000000;
filter4[42][1][1] = 35'b00000101101010101011101100010000000;
filter4[42][1][2] = 35'b11111100001101101110011100101100000;
filter4[42][2][0] = 35'b11111011011110011111000111110000000;
filter4[42][2][1] = 35'b00000000010001111001001001001000100;
filter4[42][2][2] = 35'b00001001110111100100000100100000000;
filter4[43][0][0] = 35'b00000110000111001111011110010000000;
filter4[43][0][1] = 35'b11111111001100111011010001101000000;
filter4[43][0][2] = 35'b11111111111001000011111011011101010;
filter4[43][1][0] = 35'b00000011101000111011110010110100000;
filter4[43][1][1] = 35'b00001101010101111100010101110000000;
filter4[43][1][2] = 35'b00000001100100110000100001010000000;
filter4[43][2][0] = 35'b00000011100010111110001010000000000;
filter4[43][2][1] = 35'b00001100110010011010010010100000000;
filter4[43][2][2] = 35'b11111001101001000110101100010000000;
filter4[44][0][0] = 35'b00000010010010000011101101001100000;
filter4[44][0][1] = 35'b00000101011011010000000100000000000;
filter4[44][0][2] = 35'b00000010101010010000101001010000000;
filter4[44][1][0] = 35'b11111011100011101101000011111000000;
filter4[44][1][1] = 35'b11111110011110000001100001100010000;
filter4[44][1][2] = 35'b11110101001100001001011001000000000;
filter4[44][2][0] = 35'b11111011001001000110001111011000000;
filter4[44][2][1] = 35'b11111110000001100001011100100000000;
filter4[44][2][2] = 35'b11111111000011000010001101001000000;
filter4[45][0][0] = 35'b00001000100111011100000010000000000;
filter4[45][0][1] = 35'b00000001001010001111101111011000000;
filter4[45][0][2] = 35'b11110111000100101000000010010000000;
filter4[45][1][0] = 35'b00000010111010111100111100101100000;
filter4[45][1][1] = 35'b00001111101110011000101111010000000;
filter4[45][1][2] = 35'b00000010100101110101010101010100000;
filter4[45][2][0] = 35'b00000101101010111010110010111000000;
filter4[45][2][1] = 35'b00000110100010010010101000111000000;
filter4[45][2][2] = 35'b00000011001110111100100110100000000;
filter4[46][0][0] = 35'b11111101101110100101101011100000000;
filter4[46][0][1] = 35'b11111100011000000101110100110100000;
filter4[46][0][2] = 35'b11111010001011111111111100010000000;
filter4[46][1][0] = 35'b00000000010101000110100101000010000;
filter4[46][1][1] = 35'b11111110001101111011010110010010000;
filter4[46][1][2] = 35'b11111100100011000101001000111100000;
filter4[46][2][0] = 35'b11111100110000111011011110011000000;
filter4[46][2][1] = 35'b00000111011111100011101111101000000;
filter4[46][2][2] = 35'b00000000111001000001000111100010000;
filter4[47][0][0] = 35'b00000001010111100110111011010110000;
filter4[47][0][1] = 35'b11111010100000011101110110100000000;
filter4[47][0][2] = 35'b11111011111010111110011010011000000;
filter4[47][1][0] = 35'b00001010110111010101000101100000000;
filter4[47][1][1] = 35'b00000101010110001101010000101000000;
filter4[47][1][2] = 35'b11111110100010001011001001111000000;
filter4[47][2][0] = 35'b11111111111111000110111111101000001;
filter4[47][2][1] = 35'b00001110010110111000001001000000000;
filter4[47][2][2] = 35'b11111101011011001111011100000100000;
filter4[48][0][0] = 35'b00000101000001101111011010000000000;
filter4[48][0][1] = 35'b11110110000100010000111011010000000;
filter4[48][0][2] = 35'b00000101100011010100100110110000000;
filter4[48][1][0] = 35'b00000000010111111101101101000011100;
filter4[48][1][1] = 35'b11110010111111000101101101010000000;
filter4[48][1][2] = 35'b00000010101001011111111000100000000;
filter4[48][2][0] = 35'b00000010111100000010000100001000000;
filter4[48][2][1] = 35'b11111110110000000110100001011110000;
filter4[48][2][2] = 35'b11111101101101010011011101111000000;
filter4[49][0][0] = 35'b00000001011000001101101100000110000;
filter4[49][0][1] = 35'b11111100000000111100000001101100000;
filter4[49][0][2] = 35'b11111011011111011111001100011000000;
filter4[49][1][0] = 35'b11110000100111111001010111100000000;
filter4[49][1][1] = 35'b11110110110011100010001001100000000;
filter4[49][1][2] = 35'b00000010101000000101111111100000000;
filter4[49][2][0] = 35'b00000100101000000100010010110000000;
filter4[49][2][1] = 35'b00000110100001001110011111001000000;
filter4[49][2][2] = 35'b11111101000101011001101110111100000;
filter4[50][0][0] = 35'b00000000010001100011101010100010000;
filter4[50][0][1] = 35'b11111110000000100011000111000100000;
filter4[50][0][2] = 35'b00000111001110111011011011010000000;
filter4[50][1][0] = 35'b00001001110100110000111111100000000;
filter4[50][1][1] = 35'b00001001110101111100011011100000000;
filter4[50][1][2] = 35'b11111010101011111110110111111000000;
filter4[50][2][0] = 35'b00001010001110101101001101110000000;
filter4[50][2][1] = 35'b00000100010001100100010110100000000;
filter4[50][2][2] = 35'b00001000001000110111111000000000000;
filter4[51][0][0] = 35'b00000001101101111110011001100010000;
filter4[51][0][1] = 35'b11111101111110010101001111110100000;
filter4[51][0][2] = 35'b00000111000001000111100111011000000;
filter4[51][1][0] = 35'b11110110010111100000000111010000000;
filter4[51][1][1] = 35'b11110010010011010001100010010000000;
filter4[51][1][2] = 35'b00000001001011011110100011100010000;
filter4[51][2][0] = 35'b11111011000001010001010110110000000;
filter4[51][2][1] = 35'b11111111000110101000000100011111000;
filter4[51][2][2] = 35'b11111011011001101001111001000000000;
filter4[52][0][0] = 35'b00000010101000010110111110110100000;
filter4[52][0][1] = 35'b00000110101000111010001001001000000;
filter4[52][0][2] = 35'b00000101001010001110110110100000000;
filter4[52][1][0] = 35'b11111100111110010110011101100100000;
filter4[52][1][1] = 35'b00000011001000001110111111100100000;
filter4[52][1][2] = 35'b11111110100101000000000000100000000;
filter4[52][2][0] = 35'b00001001010001110100110011010000000;
filter4[52][2][1] = 35'b11111111110101101110001010000001000;
filter4[52][2][2] = 35'b00000011000001111011111110101100000;
filter4[53][0][0] = 35'b11111001111001100101111010111000000;
filter4[53][0][1] = 35'b00000001101001100100010011100000000;
filter4[53][0][2] = 35'b11110111001010010100000001100000000;
filter4[53][1][0] = 35'b11110101010001000111010110110000000;
filter4[53][1][1] = 35'b11110011001110011001100111100000000;
filter4[53][1][2] = 35'b11110101101000110101111110100000000;
filter4[53][2][0] = 35'b00000000011111010111010111101010000;
filter4[53][2][1] = 35'b11111111101010100100011001000000100;
filter4[53][2][2] = 35'b11111111000000110000110111101111000;
filter4[54][0][0] = 35'b00000011000110000110110010100000000;
filter4[54][0][1] = 35'b11111100110001100011011100100000000;
filter4[54][0][2] = 35'b11111001010100100100000110000000000;
filter4[54][1][0] = 35'b00001000111111000000000111010000000;
filter4[54][1][1] = 35'b11111101010100010111001101110000000;
filter4[54][1][2] = 35'b00000010000011110000111100011000000;
filter4[54][2][0] = 35'b00001000100101000101000100010000000;
filter4[54][2][1] = 35'b00000110001111110000011100000000000;
filter4[54][2][2] = 35'b11111101111001011000000010011000000;
filter4[55][0][0] = 35'b00000101000101111110101101111000000;
filter4[55][0][1] = 35'b11111001011111101001111111101000000;
filter4[55][0][2] = 35'b00000001111101001110110010100100000;
filter4[55][1][0] = 35'b11111100000000111111100110011100000;
filter4[55][1][1] = 35'b11110100010000001001011100010000000;
filter4[55][1][2] = 35'b00000011111111000001001000001100000;
filter4[55][2][0] = 35'b00000000111001010000111110101100000;
filter4[55][2][1] = 35'b00000001110010100101000001110110000;
filter4[55][2][2] = 35'b11111101010101111001010001000000000;
filter4[56][0][0] = 35'b00000100110011111001001001101000000;
filter4[56][0][1] = 35'b00000000101110010001000100011100000;
filter4[56][0][2] = 35'b00000111001111101000011000101000000;
filter4[56][1][0] = 35'b00000101001101100010001100010000000;
filter4[56][1][1] = 35'b11111011100101110000100111010000000;
filter4[56][1][2] = 35'b00000010111101010001011010110000000;
filter4[56][2][0] = 35'b11111001101010101111001011111000000;
filter4[56][2][1] = 35'b11111000001110111010000011011000000;
filter4[56][2][2] = 35'b11110111101100100111001111110000000;
filter4[57][0][0] = 35'b00000011000110111100001011110000000;
filter4[57][0][1] = 35'b00000101111011111111101101111000000;
filter4[57][0][2] = 35'b00000010001000110011010101111000000;
filter4[57][1][0] = 35'b00000110000101010100110000110000000;
filter4[57][1][1] = 35'b00000111011011101101000111000000000;
filter4[57][1][2] = 35'b11111000011001111111111101011000000;
filter4[57][2][0] = 35'b11111010111010001111111110000000000;
filter4[57][2][1] = 35'b11110011010011110000100101000000000;
filter4[57][2][2] = 35'b00000001100101000011101110111100000;
filter4[58][0][0] = 35'b00000011110010101001011100100000000;
filter4[58][0][1] = 35'b11111011100111011011101111111000000;
filter4[58][0][2] = 35'b11111100110110011000101000111100000;
filter4[58][1][0] = 35'b00000001100001001000111001011010000;
filter4[58][1][1] = 35'b11111111111010011010000110011110011;
filter4[58][1][2] = 35'b11111111001101011001110111110111000;
filter4[58][2][0] = 35'b11111110100111101011110101110010000;
filter4[58][2][1] = 35'b11111101100011000000100010100000000;
filter4[58][2][2] = 35'b00000000011101000101101100110000000;
filter4[59][0][0] = 35'b11111111010011010110001000101111000;
filter4[59][0][1] = 35'b00000010011111111110011001010000000;
filter4[59][0][2] = 35'b00000100011100111101110000100000000;
filter4[59][1][0] = 35'b00000111001111000101111001000000000;
filter4[59][1][1] = 35'b00000010101101011001110111110100000;
filter4[59][1][2] = 35'b11111010111111110111100111001000000;
filter4[59][2][0] = 35'b11111000110110011100001001110000000;
filter4[59][2][1] = 35'b11110010010001011011101110100000000;
filter4[59][2][2] = 35'b11111010000101110101100001010000000;
filter4[60][0][0] = 35'b11111111111111010010111101100100010;
filter4[60][0][1] = 35'b11111110001011110010000101101010000;
filter4[60][0][2] = 35'b11111100111110110010100101001100000;
filter4[60][1][0] = 35'b00000000000100110011000110101010111;
filter4[60][1][1] = 35'b11111110111100000101101100010100000;
filter4[60][1][2] = 35'b11111110010101011010100001011000000;
filter4[60][2][0] = 35'b11111110101011100101011110110000000;
filter4[60][2][1] = 35'b11111110110010001011100101000110000;
filter4[60][2][2] = 35'b11111110000110011101001100111100000;
filter4[61][0][0] = 35'b00000001100011111101000100101010000;
filter4[61][0][1] = 35'b00001000001011101001001101010000000;
filter4[61][0][2] = 35'b11111110110001011101010001010010000;
filter4[61][1][0] = 35'b00001001010011111110011110100000000;
filter4[61][1][1] = 35'b00000011101001000110101011111000000;
filter4[61][1][2] = 35'b11111011111110111111010101000000000;
filter4[61][2][0] = 35'b00000010100101011101101101011000000;
filter4[61][2][1] = 35'b11111010101010011100111111111000000;
filter4[61][2][2] = 35'b11111011001100011010001011001000000;
filter4[62][0][0] = 35'b11111110110001010111001100011100000;
filter4[62][0][1] = 35'b00000000001110001100100000110100010;
filter4[62][0][2] = 35'b00000100101011110111001010111000000;
filter4[62][1][0] = 35'b00000001011100100111001101011000000;
filter4[62][1][1] = 35'b00000000000011001111110010111000110;
filter4[62][1][2] = 35'b00000000010011000100010111000011000;
filter4[62][2][0] = 35'b00000101010011110110101011001000000;
filter4[62][2][1] = 35'b11111110010010010000000100000010000;
filter4[62][2][2] = 35'b11111000100111010001001101001000000;
filter4[63][0][0] = 35'b00000011101011000100011000101100000;
filter4[63][0][1] = 35'b00000111101011101110100011100000000;
filter4[63][0][2] = 35'b00001001011111101000011100100000000;
filter4[63][1][0] = 35'b00000010111010100110100001110100000;
filter4[63][1][1] = 35'b11111100100110110001011001011100000;
filter4[63][1][2] = 35'b00000100011000010101111100111000000;
filter4[63][2][0] = 35'b11111100010100101010001101101100000;
filter4[63][2][1] = 35'b11110111100110001101100011010000000;
filter4[63][2][2] = 35'b11110011101011110101010110100000000;
filter4[64][0][0] = 35'b00000000000011001101000001011101000;
filter4[64][0][1] = 35'b00000110101101011001111011100000000;
filter4[64][0][2] = 35'b11111100111101101011000001111100000;
filter4[64][1][0] = 35'b00000000000001001110100001001110000;
filter4[64][1][1] = 35'b11111111010011011010111001010100000;
filter4[64][1][2] = 35'b11110100101010011000010010110000000;
filter4[64][2][0] = 35'b00000101110010111110111001010000000;
filter4[64][2][1] = 35'b11111110011101101001100000111010000;
filter4[64][2][2] = 35'b11111111000110001001110100110110000;
filter4[65][0][0] = 35'b00000010000011011011110101101000000;
filter4[65][0][1] = 35'b00000100100100000100101110001000000;
filter4[65][0][2] = 35'b11111100100001010011010010110100000;
filter4[65][1][0] = 35'b11111111101000110100011011101111000;
filter4[65][1][1] = 35'b00000010100101011011111011010000000;
filter4[65][1][2] = 35'b11111100011100110000101100100100000;
filter4[65][2][0] = 35'b00000000100111001010101000111011000;
filter4[65][2][1] = 35'b00000110100101110110100111110000000;
filter4[65][2][2] = 35'b11111011100110000010101110010000000;
filter4[66][0][0] = 35'b11111111011110100010111111111000000;
filter4[66][0][1] = 35'b11110100101000011011100000010000000;
filter4[66][0][2] = 35'b00000110010110000101010100001000000;
filter4[66][1][0] = 35'b00000001100000001110000101011110000;
filter4[66][1][1] = 35'b11111101001010111111000001100100000;
filter4[66][1][2] = 35'b11111110110000010011011101100000000;
filter4[66][2][0] = 35'b11111111110011111011011000001110100;
filter4[66][2][1] = 35'b00010000111010111100011110000000000;
filter4[66][2][2] = 35'b00000011111111101011010010001000000;
filter4[67][0][0] = 35'b11111110010100001100110001010110000;
filter4[67][0][1] = 35'b00001011000000101111000011100000000;
filter4[67][0][2] = 35'b11111001110001010001110101111000000;
filter4[67][1][0] = 35'b11111101011110011100100110001000000;
filter4[67][1][1] = 35'b00000100011011010010000110011000000;
filter4[67][1][2] = 35'b11111010001010110101101111011000000;
filter4[67][2][0] = 35'b00000101010010100101110111100000000;
filter4[67][2][1] = 35'b11111111001010110111111001111000000;
filter4[67][2][2] = 35'b11111101011000100111101100000100000;
filter4[68][0][0] = 35'b11111011000010101101101001100000000;
filter4[68][0][1] = 35'b00000011111111100100101000110100000;
filter4[68][0][2] = 35'b00000100110001001000001001101000000;
filter4[68][1][0] = 35'b11111101100001010111011001100000000;
filter4[68][1][1] = 35'b00000010011110110010001110000100000;
filter4[68][1][2] = 35'b00000001000100000100110111111000000;
filter4[68][2][0] = 35'b00000100001111111000110011000000000;
filter4[68][2][1] = 35'b11111010100100100000101111011000000;
filter4[68][2][2] = 35'b11111110111010011010110110100110000;
filter4[69][0][0] = 35'b11111010000101000111111000010000000;
filter4[69][0][1] = 35'b00000000001001010110100111001011110;
filter4[69][0][2] = 35'b00000010111010000011101000111000000;
filter4[69][1][0] = 35'b11111100010000110100111011100100000;
filter4[69][1][1] = 35'b00000001110101011011000111110100000;
filter4[69][1][2] = 35'b00000011100000110111110001101100000;
filter4[69][2][0] = 35'b11111111010000011110110011101010000;
filter4[69][2][1] = 35'b00000011010000010110010001111100000;
filter4[69][2][2] = 35'b11111111010110000111100100111101000;
filter4[70][0][0] = 35'b11111000101111000000111100100000000;
filter4[70][0][1] = 35'b00000000110000111100111010000010000;
filter4[70][0][2] = 35'b00001000110101100110001110100000000;
filter4[70][1][0] = 35'b11111001010000111101010111101000000;
filter4[70][1][1] = 35'b00000101101011011011110001001000000;
filter4[70][1][2] = 35'b00000111010110011001111111010000000;
filter4[70][2][0] = 35'b11111011110011110111001001101000000;
filter4[70][2][1] = 35'b00000011101010010111011100100100000;
filter4[70][2][2] = 35'b00000011100000111100111101110100000;
filter4[71][0][0] = 35'b00000000111100010001001100110010000;
filter4[71][0][1] = 35'b00001000111110011100011000010000000;
filter4[71][0][2] = 35'b11110110111000110111100000010000000;
filter4[71][1][0] = 35'b11111100000011101011110011011100000;
filter4[71][1][1] = 35'b00000010100010010001101101110000000;
filter4[71][1][2] = 35'b11111001111010010010111000011000000;
filter4[71][2][0] = 35'b00000011111011010000000110100000000;
filter4[71][2][1] = 35'b11111101010001010001011011000000000;
filter4[71][2][2] = 35'b11111111011110101111011011111111000;
filter4[72][0][0] = 35'b00000001011100111101010011111100000;
filter4[72][0][1] = 35'b11111100101110100001000011110100000;
filter4[72][0][2] = 35'b00000111010101001011001001111000000;
filter4[72][1][0] = 35'b00000111111000110101010101010000000;
filter4[72][1][1] = 35'b00000001000010100001110111000100000;
filter4[72][1][2] = 35'b11111011111011100110010111101000000;
filter4[72][2][0] = 35'b00000101100001101010000000100000000;
filter4[72][2][1] = 35'b11111110011111100010000001000000000;
filter4[72][2][2] = 35'b11111000110000100111111010111000000;
filter4[73][0][0] = 35'b00001000110101111001000101100000000;
filter4[73][0][1] = 35'b00000000111110000110101100001111000;
filter4[73][0][2] = 35'b00000110001111010100110000010000000;
filter4[73][1][0] = 35'b11111111110010111010011011111001010;
filter4[73][1][1] = 35'b11111111000010111100111111110000000;
filter4[73][1][2] = 35'b00000011110000000111111111111100000;
filter4[73][2][0] = 35'b00000000010000100010110001011100000;
filter4[73][2][1] = 35'b11111111111001001111101000000011000;
filter4[73][2][2] = 35'b11110110101101110010010010010000000;
filter4[74][0][0] = 35'b11111100100100111011000101000100000;
filter4[74][0][1] = 35'b11111111000011100111000110111110000;
filter4[74][0][2] = 35'b11111000010010110011101011011000000;
filter4[74][1][0] = 35'b11111001110111010101110101110000000;
filter4[74][1][1] = 35'b11111001001110000000100011100000000;
filter4[74][1][2] = 35'b11110101100010111000010101010000000;
filter4[74][2][0] = 35'b00000111010100110110110110101000000;
filter4[74][2][1] = 35'b00000110000011111000001010101000000;
filter4[74][2][2] = 35'b00001000110011010101111010010000000;
filter4[75][0][0] = 35'b00000110111110111110111011101000000;
filter4[75][0][1] = 35'b00000111110011010101101100101000000;
filter4[75][0][2] = 35'b00000110010101000110001010001000000;
filter4[75][1][0] = 35'b00000101111011110001000111101000000;
filter4[75][1][1] = 35'b11111101111101111010001101000100000;
filter4[75][1][2] = 35'b11111101001100110100010010111000000;
filter4[75][2][0] = 35'b00000010011001100001100011100000000;
filter4[75][2][1] = 35'b11111111000000010111100010111101000;
filter4[75][2][2] = 35'b11110100010000100001001011000000000;
filter4[76][0][0] = 35'b11111001001001001110011101100000000;
filter4[76][0][1] = 35'b11111011110111101100111111101000000;
filter4[76][0][2] = 35'b11111100111101001000100011000000000;
filter4[76][1][0] = 35'b00000000001010001011000101111000010;
filter4[76][1][1] = 35'b11111100110101100001000101010100000;
filter4[76][1][2] = 35'b00000000111010101101000011100000000;
filter4[76][2][0] = 35'b00000011001101101100010000000000000;
filter4[76][2][1] = 35'b11111010000011101011101000001000000;
filter4[76][2][2] = 35'b11111110011101001101000111000110000;
filter4[77][0][0] = 35'b00000010011101111010010110100000000;
filter4[77][0][1] = 35'b11111111100011101000100010111001100;
filter4[77][0][2] = 35'b00000000111111011011110001110001000;
filter4[77][1][0] = 35'b00000011001100000010000011111000000;
filter4[77][1][1] = 35'b00000000101001101001000010110011000;
filter4[77][1][2] = 35'b11111111001000111100101101000111000;
filter4[77][2][0] = 35'b00001001100010111001100000100000000;
filter4[77][2][1] = 35'b00000010111111001000011010011000000;
filter4[77][2][2] = 35'b11111010101110111000101110011000000;
filter4[78][0][0] = 35'b11111110100000000101111001011010000;
filter4[78][0][1] = 35'b11111001101001000001110011001000000;
filter4[78][0][2] = 35'b11111000010101110011110110011000000;
filter4[78][1][0] = 35'b11111110010000011101011111101110000;
filter4[78][1][1] = 35'b11111100010000110111101000101100000;
filter4[78][1][2] = 35'b00000001011110011011110010100100000;
filter4[78][2][0] = 35'b00000111100010100100111000111000000;
filter4[78][2][1] = 35'b00000010111101011000110111110100000;
filter4[78][2][2] = 35'b00000001010001011110011001000110000;
filter4[79][0][0] = 35'b11111011110000110110010101011000000;
filter4[79][0][1] = 35'b00000001011101011000011000110010000;
filter4[79][0][2] = 35'b00000111110111010111101100110000000;
filter4[79][1][0] = 35'b00000011001110001011010011100100000;
filter4[79][1][1] = 35'b00000011001010100100100110111000000;
filter4[79][1][2] = 35'b11111100101011111011111110011000000;
filter4[79][2][0] = 35'b00000000101111110100010001100101000;
filter4[79][2][1] = 35'b11111100010111111110011101100100000;
filter4[79][2][2] = 35'b11110101100001011100111110100000000;
filter4[80][0][0] = 35'b00000010010010101100010110101100000;
filter4[80][0][1] = 35'b00000011101110000000010111100000000;
filter4[80][0][2] = 35'b11111111111001000110100110100000110;
filter4[80][1][0] = 35'b11111111100100000011010111011101100;
filter4[80][1][1] = 35'b00000101001011001010011111101000000;
filter4[80][1][2] = 35'b11111100011100100110010010001000000;
filter4[80][2][0] = 35'b00000011111010010011111111010000000;
filter4[80][2][1] = 35'b11111101000110101001000111011100000;
filter4[80][2][2] = 35'b11110011100001111011011110000000000;
filter4[81][0][0] = 35'b11111111011001111010010010101010000;
filter4[81][0][1] = 35'b00000000100101111001001010000010000;
filter4[81][0][2] = 35'b00000001101100110001101000110100000;
filter4[81][1][0] = 35'b11111111100101101010000010111011000;
filter4[81][1][1] = 35'b00000000101111100101101010111111000;
filter4[81][1][2] = 35'b11111011100111011111111100100000000;
filter4[81][2][0] = 35'b00000100001111000000000110001000000;
filter4[81][2][1] = 35'b00000110101100000000110111010000000;
filter4[81][2][2] = 35'b11111000011011011000001010001000000;
filter4[82][0][0] = 35'b00000110110010101001010011011000000;
filter4[82][0][1] = 35'b00000101001001011111001011101000000;
filter4[82][0][2] = 35'b00000001110011001001001011111110000;
filter4[82][1][0] = 35'b00000110101011101101111001001000000;
filter4[82][1][1] = 35'b00000110011000011100011010101000000;
filter4[82][1][2] = 35'b00000011000101010111001010110100000;
filter4[82][2][0] = 35'b11111111001100100110111100000001000;
filter4[82][2][1] = 35'b00000000101100110000001111010110000;
filter4[82][2][2] = 35'b00000000000101101011000111000100101;
filter4[83][0][0] = 35'b11111011100000110011001010000000000;
filter4[83][0][1] = 35'b00000101011000000110110110110000000;
filter4[83][0][2] = 35'b00000011000100111101000011110100000;
filter4[83][1][0] = 35'b11111100111101011010000000010100000;
filter4[83][1][1] = 35'b11111101000010110001011111011100000;
filter4[83][1][2] = 35'b11111001111011000100011101101000000;
filter4[83][2][0] = 35'b11111110011111110101000010110100000;
filter4[83][2][1] = 35'b00000111100101111111000000110000000;
filter4[83][2][2] = 35'b11110110101011011011110011110000000;
filter4[84][0][0] = 35'b00000011110001010000010111010100000;
filter4[84][0][1] = 35'b00000000101011001010000001101010000;
filter4[84][0][2] = 35'b00000000101010100001100001000110000;
filter4[84][1][0] = 35'b00000010111011111001111110100100000;
filter4[84][1][1] = 35'b00001000001110011100100001000000000;
filter4[84][1][2] = 35'b00000001010000010000110111001110000;
filter4[84][2][0] = 35'b00000010011011100011110100100000000;
filter4[84][2][1] = 35'b11111111001101000001100001110011000;
filter4[84][2][2] = 35'b00000000101101110000101111100010000;
filter4[85][0][0] = 35'b11111001010001101101001011011000000;
filter4[85][0][1] = 35'b00000100111111010010010010010000000;
filter4[85][0][2] = 35'b00000101011111010010110101000000000;
filter4[85][1][0] = 35'b00000100011110011010001111001000000;
filter4[85][1][1] = 35'b11111101001110010011010111001000000;
filter4[85][1][2] = 35'b00000010000111100011110101001100000;
filter4[85][2][0] = 35'b11111110010110011110000111111010000;
filter4[85][2][1] = 35'b00001000101010011111011110110000000;
filter4[85][2][2] = 35'b11111111000001111101001110110100000;
filter4[86][0][0] = 35'b00000010111110001000100000110100000;
filter4[86][0][1] = 35'b00000101101100101001110100100000000;
filter4[86][0][2] = 35'b00000011100110110100000101001000000;
filter4[86][1][0] = 35'b11111101101100111011011010101000000;
filter4[86][1][1] = 35'b00000000011000000010011010001111100;
filter4[86][1][2] = 35'b00000010101110110000011011111100000;
filter4[86][2][0] = 35'b00000111001100111010001001100000000;
filter4[86][2][1] = 35'b00000010010001001011000111111100000;
filter4[86][2][2] = 35'b11111111000110000101011111000111000;
filter4[87][0][0] = 35'b11111110011110100000011100100100000;
filter4[87][0][1] = 35'b00000001110011101100001101010000000;
filter4[87][0][2] = 35'b00000100011001001000111111011000000;
filter4[87][1][0] = 35'b11111011001100100011101001101000000;
filter4[87][1][1] = 35'b00000000110111100010110111100101000;
filter4[87][1][2] = 35'b11111011100100001111101010110000000;
filter4[87][2][0] = 35'b00000100011110100110001001101000000;
filter4[87][2][1] = 35'b11111101111110101110111000011100000;
filter4[87][2][2] = 35'b11110001001111101100111011110000000;
filter4[88][0][0] = 35'b00001001110001001101000100110000000;
filter4[88][0][1] = 35'b00000010010010110000011110110100000;
filter4[88][0][2] = 35'b11111101011011011000101000110000000;
filter4[88][1][0] = 35'b00000100011110110010111011100000000;
filter4[88][1][1] = 35'b00000010110111010111101110011000000;
filter4[88][1][2] = 35'b11111111001011111001111011110100000;
filter4[88][2][0] = 35'b11111111010001000101111010010111000;
filter4[88][2][1] = 35'b00000101011101101110110000010000000;
filter4[88][2][2] = 35'b11111101110100010001010110101000000;
filter4[89][0][0] = 35'b00000101000001110010000100010000000;
filter4[89][0][1] = 35'b00000011110111100110001000011000000;
filter4[89][0][2] = 35'b00000011000111010000111011010100000;
filter4[89][1][0] = 35'b00000100111111111001010001110000000;
filter4[89][1][1] = 35'b00000100010001111100110010000000000;
filter4[89][1][2] = 35'b00000100010011000101100110110000000;
filter4[89][2][0] = 35'b11111011110100011011111110111000000;
filter4[89][2][1] = 35'b00000110000010110111001000000000000;
filter4[89][2][2] = 35'b00000010001001101110000111100000000;
filter4[90][0][0] = 35'b11111101101000111000111011110100000;
filter4[90][0][1] = 35'b00000001011000110111110101010010000;
filter4[90][0][2] = 35'b11111010101101000011010110000000000;
filter4[90][1][0] = 35'b11111110110011000001001100010010000;
filter4[90][1][1] = 35'b11111011001110000010100101100000000;
filter4[90][1][2] = 35'b11111000100100011111101001100000000;
filter4[90][2][0] = 35'b00000100011100110001001110011000000;
filter4[90][2][1] = 35'b11111000111011100011001101101000000;
filter4[90][2][2] = 35'b11111011001111001101010101110000000;
filter4[91][0][0] = 35'b00001001110001111010101000100000000;
filter4[91][0][1] = 35'b00001011000010101001110011100000000;
filter4[91][0][2] = 35'b00000010001110101001101101100100000;
filter4[91][1][0] = 35'b00000011110110101101000100111100000;
filter4[91][1][1] = 35'b00001000011101011111100000000000000;
filter4[91][1][2] = 35'b00000101101110011111101001110000000;
filter4[91][2][0] = 35'b11111110111100000111010101110000000;
filter4[91][2][1] = 35'b00001101010100100100010101100000000;
filter4[91][2][2] = 35'b00000100000110100001001010000000000;
filter4[92][0][0] = 35'b11111010011111111001001001011000000;
filter4[92][0][1] = 35'b00000111011001111110100000100000000;
filter4[92][0][2] = 35'b00000011010101001011101110110000000;
filter4[92][1][0] = 35'b11111011000100010111111000011000000;
filter4[92][1][1] = 35'b11111100010011110010110001011000000;
filter4[92][1][2] = 35'b00000110001100110100011001011000000;
filter4[92][2][0] = 35'b00000000001001111100001101000110110;
filter4[92][2][1] = 35'b11111101000011111000011110010000000;
filter4[92][2][2] = 35'b00000000111111010000110101010100000;
filter4[93][0][0] = 35'b00000100011010000001110101110000000;
filter4[93][0][1] = 35'b00010111101001100000000111100000000;
filter4[93][0][2] = 35'b11111110111111001100111000110100000;
filter4[93][1][0] = 35'b00000100001000101101000001110000000;
filter4[93][1][1] = 35'b00001011010000100110111001100000000;
filter4[93][1][2] = 35'b00000110101000011111010100011000000;
filter4[93][2][0] = 35'b11111100000010100100111000000100000;
filter4[93][2][1] = 35'b00000101110010111110000110000000000;
filter4[93][2][2] = 35'b00001110101011001100001100110000000;
filter4[94][0][0] = 35'b11111110110111101011111001001110000;
filter4[94][0][1] = 35'b11111011101111010101011001110000000;
filter4[94][0][2] = 35'b11111100110111110001101101110100000;
filter4[94][1][0] = 35'b00000101011111110010111100000000000;
filter4[94][1][1] = 35'b00000101110000000010000111111000000;
filter4[94][1][2] = 35'b11111011100001101100111111011000000;
filter4[94][2][0] = 35'b11111101111010101010011000000100000;
filter4[94][2][1] = 35'b11111111110001110010111101001110110;
filter4[94][2][2] = 35'b11111111101100101101001110111010000;
filter4[95][0][0] = 35'b00001111000010101100111010000000000;
filter4[95][0][1] = 35'b11111111010100110110000100001001000;
filter4[95][0][2] = 35'b00000100101001010110100101110000000;
filter4[95][1][0] = 35'b00000010100010111111011100010100000;
filter4[95][1][1] = 35'b00000001111111101101001010101000000;
filter4[95][1][2] = 35'b11111010100101000101000011011000000;
filter4[95][2][0] = 35'b11111101110111001100100100110000000;
filter4[95][2][1] = 35'b00010011001001001000011010100000000;
filter4[95][2][2] = 35'b00000011001001010101000110111100000;
filter4[96][0][0] = 35'b00000010000100110111001110010100000;
filter4[96][0][1] = 35'b00000000001000101001000000101100110;
filter4[96][0][2] = 35'b11111011110100111011110100110000000;
filter4[96][1][0] = 35'b11111101101001101101010100100100000;
filter4[96][1][1] = 35'b11110101011111000100111110110000000;
filter4[96][1][2] = 35'b11111111101110001001011100111010000;
filter4[96][2][0] = 35'b11111000000110000000101101110000000;
filter4[96][2][1] = 35'b11111100101000000011010100100000000;
filter4[96][2][2] = 35'b00001010001000111110111101000000000;
filter4[97][0][0] = 35'b00000100010001101011100101110000000;
filter4[97][0][1] = 35'b11111111010001010110001110101001000;
filter4[97][0][2] = 35'b11111101110101000010100000110100000;
filter4[97][1][0] = 35'b00000010111101001011111011010000000;
filter4[97][1][1] = 35'b11111011110100000101011000010000000;
filter4[97][1][2] = 35'b11111100001010100000001100000000000;
filter4[97][2][0] = 35'b11111011100010001010000010001000000;
filter4[97][2][1] = 35'b11111100100101111100001011101000000;
filter4[97][2][2] = 35'b00000110001110010001010100010000000;
filter4[98][0][0] = 35'b00000010010010111011001110101000000;
filter4[98][0][1] = 35'b11110111011111111100110000100000000;
filter4[98][0][2] = 35'b11111100000001110100000000111100000;
filter4[98][1][0] = 35'b00000001111001001110111010010100000;
filter4[98][1][1] = 35'b11111100110000100011111010010000000;
filter4[98][1][2] = 35'b00000100111110001100110001100000000;
filter4[98][2][0] = 35'b11111000101110000100100110101000000;
filter4[98][2][1] = 35'b00000000111001111111000100101100000;
filter4[98][2][2] = 35'b00000110010100011010000001011000000;
filter4[99][0][0] = 35'b00000110000010110010101001110000000;
filter4[99][0][1] = 35'b00000010000011000110100111001100000;
filter4[99][0][2] = 35'b11111001100101100110100100101000000;
filter4[99][1][0] = 35'b00000001010011000010100110100110000;
filter4[99][1][1] = 35'b11110101110101101000010001110000000;
filter4[99][1][2] = 35'b11111100010010101011001111100100000;
filter4[99][2][0] = 35'b11111010011101111011110101000000000;
filter4[99][2][1] = 35'b11111101101011100110111111011000000;
filter4[99][2][2] = 35'b00001001010101010010001000000000000;
filter4[100][0][0] = 35'b00000101000001001011011010011000000;
filter4[100][0][1] = 35'b11111101001100001001110111111100000;
filter4[100][0][2] = 35'b00000011111111101001111101000000000;
filter4[100][1][0] = 35'b11111001110111001101100100000000000;
filter4[100][1][1] = 35'b11111111101111001101011001010010000;
filter4[100][1][2] = 35'b11111111100110000000110010100101000;
filter4[100][2][0] = 35'b11111110110111101001000101001000000;
filter4[100][2][1] = 35'b00000100001000101110000000000000000;
filter4[100][2][2] = 35'b00000001010100010011001100101110000;
filter4[101][0][0] = 35'b00000111100100110011111110000000000;
filter4[101][0][1] = 35'b00000100110000010111001011110000000;
filter4[101][0][2] = 35'b11111110010011010001010001011000000;
filter4[101][1][0] = 35'b00001100011010101101100001110000000;
filter4[101][1][1] = 35'b11111111110000100111110110111000100;
filter4[101][1][2] = 35'b11111001010110010110111100110000000;
filter4[101][2][0] = 35'b00000100000100111111111011100000000;
filter4[101][2][1] = 35'b11111010001001100110110000000000000;
filter4[101][2][2] = 35'b00000011100000100000010011110100000;
filter4[102][0][0] = 35'b11111110000110001001100101101000000;
filter4[102][0][1] = 35'b00001101011110010111110010000000000;
filter4[102][0][2] = 35'b00000100101101111110101010001000000;
filter4[102][1][0] = 35'b00000010111010110001110010001100000;
filter4[102][1][1] = 35'b00000101110001011100101101111000000;
filter4[102][1][2] = 35'b00000001111100100101111001001000000;
filter4[102][2][0] = 35'b00000010001100000111000000110000000;
filter4[102][2][1] = 35'b00000001010000100111001011110110000;
filter4[102][2][2] = 35'b00000011100100001011110110010000000;
filter4[103][0][0] = 35'b00000011000011000011100110101100000;
filter4[103][0][1] = 35'b11111111011101101010111100110111000;
filter4[103][0][2] = 35'b11111110011000010101101010000010000;
filter4[103][1][0] = 35'b00000001001100101011100010010000000;
filter4[103][1][1] = 35'b11110100110011100011110111000000000;
filter4[103][1][2] = 35'b11111110001101111000001101001010000;
filter4[103][2][0] = 35'b11111101010100101101101010001100000;
filter4[103][2][1] = 35'b11111110110001010100110111011110000;
filter4[103][2][2] = 35'b00000100001100001111010000000000000;
filter4[104][0][0] = 35'b00000011101101111010000100000000000;
filter4[104][0][1] = 35'b00000001001000100111000110111000000;
filter4[104][0][2] = 35'b00000010100011010000110010111100000;
filter4[104][1][0] = 35'b00000000001011110011101010010000010;
filter4[104][1][1] = 35'b00001000011110111000000101100000000;
filter4[104][1][2] = 35'b11111110010001011011111011010000000;
filter4[104][2][0] = 35'b00000010101010010001011110001100000;
filter4[104][2][1] = 35'b11111101000111000101001111111100000;
filter4[104][2][2] = 35'b11111001011001101000001011110000000;
filter4[105][0][0] = 35'b00000000010010100011100010111010100;
filter4[105][0][1] = 35'b00000001010111011000111001111010000;
filter4[105][0][2] = 35'b00001100001010011010010110100000000;
filter4[105][1][0] = 35'b00001001010000011111000010000000000;
filter4[105][1][1] = 35'b00000111101100011001000011011000000;
filter4[105][1][2] = 35'b00000100110101101011010001101000000;
filter4[105][2][0] = 35'b00000010001000000000000110101100000;
filter4[105][2][1] = 35'b11111011110010011011111001110000000;
filter4[105][2][2] = 35'b00000011100000001000101101011000000;
filter4[106][0][0] = 35'b00000111010001011011110001010000000;
filter4[106][0][1] = 35'b00000000101100001110110100011000000;
filter4[106][0][2] = 35'b11111101010000000111010111110000000;
filter4[106][1][0] = 35'b11111000001111101100101101000000000;
filter4[106][1][1] = 35'b11111101000101110100011011010100000;
filter4[106][1][2] = 35'b11110010100011010111110110110000000;
filter4[106][2][0] = 35'b11111000011101100101000111011000000;
filter4[106][2][1] = 35'b11111001101110101101000101010000000;
filter4[106][2][2] = 35'b11110111000111110110000100010000000;
filter4[107][0][0] = 35'b00000010100011000101101001010100000;
filter4[107][0][1] = 35'b00000101100110111110010010001000000;
filter4[107][0][2] = 35'b00001101110011011111010010100000000;
filter4[107][1][0] = 35'b00000100011111110111011001100000000;
filter4[107][1][1] = 35'b00001000001000101000110000100000000;
filter4[107][1][2] = 35'b00001001101100101101110110100000000;
filter4[107][2][0] = 35'b11111111101010001110100001110100100;
filter4[107][2][1] = 35'b11111101001101100110110111001100000;
filter4[107][2][2] = 35'b00000100001111111111111110000000000;
filter4[108][0][0] = 35'b00000001111110011000111100001000000;
filter4[108][0][1] = 35'b11111110001100111101010100110100000;
filter4[108][0][2] = 35'b11111111111011010011110100111100111;
filter4[108][1][0] = 35'b11111110011101011100100010010000000;
filter4[108][1][1] = 35'b00000001110101101011110001101110000;
filter4[108][1][2] = 35'b00000011100001101111001001010100000;
filter4[108][2][0] = 35'b11111110000011101110011100010110000;
filter4[108][2][1] = 35'b00000100010000101010101111101000000;
filter4[108][2][2] = 35'b11111101010110101001011000000100000;
filter4[109][0][0] = 35'b11111100110111110100110001011000000;
filter4[109][0][1] = 35'b11111110011011011011110100011010000;
filter4[109][0][2] = 35'b00001000110100111101100101000000000;
filter4[109][1][0] = 35'b00000001100011011110001110110000000;
filter4[109][1][1] = 35'b00001000001110000001010110100000000;
filter4[109][1][2] = 35'b00000010100000000101000110110000000;
filter4[109][2][0] = 35'b00000011011110111111000011000000000;
filter4[109][2][1] = 35'b11111001111111010111011011101000000;
filter4[109][2][2] = 35'b00000101101011100101110001011000000;
filter4[110][0][0] = 35'b11111110110111101001011111000010000;
filter4[110][0][1] = 35'b11111101001011110001111000110000000;
filter4[110][0][2] = 35'b00000111011111111111011011100000000;
filter4[110][1][0] = 35'b11111101001011101000001011111000000;
filter4[110][1][1] = 35'b00000000011111011001011100100101000;
filter4[110][1][2] = 35'b11111110101010101110110000111100000;
filter4[110][2][0] = 35'b11111100010111101011001101010000000;
filter4[110][2][1] = 35'b11111110101000011011111111000110000;
filter4[110][2][2] = 35'b11111001111110000100001100110000000;
filter4[111][0][0] = 35'b11111110001000110100001111000110000;
filter4[111][0][1] = 35'b11111110000111110010010011010000000;
filter4[111][0][2] = 35'b00000110010111101110011010111000000;
filter4[111][1][0] = 35'b00000101100001000100111011011000000;
filter4[111][1][1] = 35'b00000100110100001101110101111000000;
filter4[111][1][2] = 35'b00000001010100101100111101110110000;
filter4[111][2][0] = 35'b11111110101000000100110011100010000;
filter4[111][2][1] = 35'b00000001001001100111010101110110000;
filter4[111][2][2] = 35'b11111101101000101010100010110100000;
filter4[112][0][0] = 35'b11111011101100001001010011010000000;
filter4[112][0][1] = 35'b00000010100001110011100111000000000;
filter4[112][0][2] = 35'b00000001001110100111101100011100000;
filter4[112][1][0] = 35'b11111010111000011110000101011000000;
filter4[112][1][1] = 35'b00000110001011100011001100111000000;
filter4[112][1][2] = 35'b11111101011100011111011001100000000;
filter4[112][2][0] = 35'b00000101100010110001011110100000000;
filter4[112][2][1] = 35'b00000011101110110001101000010100000;
filter4[112][2][2] = 35'b00000010101000010110111001110100000;
filter4[113][0][0] = 35'b00000110010001000110000000101000000;
filter4[113][0][1] = 35'b11111111101100000010000111011101100;
filter4[113][0][2] = 35'b00000001010011111000101111011000000;
filter4[113][1][0] = 35'b00000000010001110101000101000000100;
filter4[113][1][1] = 35'b00000110010111100010010110010000000;
filter4[113][1][2] = 35'b00001001101101011111111101110000000;
filter4[113][2][0] = 35'b00000000111001110000001000111110000;
filter4[113][2][1] = 35'b00000101010011100101110101111000000;
filter4[113][2][2] = 35'b00000111110011010010001111111000000;
filter4[114][0][0] = 35'b11110110100001111111010111010000000;
filter4[114][0][1] = 35'b11111101111001100010011111010100000;
filter4[114][0][2] = 35'b11111011010111000110000000101000000;
filter4[114][1][0] = 35'b11111010001010101110010001100000000;
filter4[114][1][1] = 35'b11111110001100111000110010011110000;
filter4[114][1][2] = 35'b11110111110010110110100000000000000;
filter4[114][2][0] = 35'b11111011011001001001000010111000000;
filter4[114][2][1] = 35'b11111010101001110011101001001000000;
filter4[114][2][2] = 35'b11111110101011000100100100111000000;
filter4[115][0][0] = 35'b11111101100000011110000010001100000;
filter4[115][0][1] = 35'b11111101111111101001011011100100000;
filter4[115][0][2] = 35'b00000100101011010101000001001000000;
filter4[115][1][0] = 35'b11111101101101010101011111001100000;
filter4[115][1][1] = 35'b00001001011010101001011100010000000;
filter4[115][1][2] = 35'b00000101110111110011100000000000000;
filter4[115][2][0] = 35'b00000000101010110010110100110110000;
filter4[115][2][1] = 35'b11111111011010111001001101101010000;
filter4[115][2][2] = 35'b00000001110110001111110000011010000;
filter4[116][0][0] = 35'b00000100110011101001011110101000000;
filter4[116][0][1] = 35'b11110100101111100111100101100000000;
filter4[116][0][2] = 35'b11111100001111111001111011111000000;
filter4[116][1][0] = 35'b11111110001001100011111110010000000;
filter4[116][1][1] = 35'b00000001010010111101110111110100000;
filter4[116][1][2] = 35'b00000001011111001001011111010110000;
filter4[116][2][0] = 35'b11111001110011100011100011010000000;
filter4[116][2][1] = 35'b11111111110011010111111010001111000;
filter4[116][2][2] = 35'b11111001101001101111111101101000000;
filter4[117][0][0] = 35'b11111110110111001111000000011110000;
filter4[117][0][1] = 35'b00000000111101101111100110010010000;
filter4[117][0][2] = 35'b11111111000111111001101000001101000;
filter4[117][1][0] = 35'b11111111110100101111010100100100110;
filter4[117][1][1] = 35'b00001000010110101101111001000000000;
filter4[117][1][2] = 35'b00000010110101110011110100100100000;
filter4[117][2][0] = 35'b11111111111100001011001101001011101;
filter4[117][2][1] = 35'b00000100101001010100110100000000000;
filter4[117][2][2] = 35'b00001000101110110111010110100000000;
filter4[118][0][0] = 35'b11110110111100011101100000100000000;
filter4[118][0][1] = 35'b11111111001100101011100010111011000;
filter4[118][0][2] = 35'b11111111011011010100101100101100000;
filter4[118][1][0] = 35'b11110110011110011101100011100000000;
filter4[118][1][1] = 35'b11111100100011111110111000111100000;
filter4[118][1][2] = 35'b11111110110010001111100011101100000;
filter4[118][2][0] = 35'b00000001101001000101100000110000000;
filter4[118][2][1] = 35'b00000111110100110010000001010000000;
filter4[118][2][2] = 35'b11111110100101010100001111110010000;
filter4[119][0][0] = 35'b11111100001010101101110001100000000;
filter4[119][0][1] = 35'b11111110001101110111110011001100000;
filter4[119][0][2] = 35'b11111111011011000001111100111010000;
filter4[119][1][0] = 35'b00000010010111010011111101010000000;
filter4[119][1][1] = 35'b00000011011001011110110010101000000;
filter4[119][1][2] = 35'b00000010110001100100111001110000000;
filter4[119][2][0] = 35'b00000001010010010101101011100010000;
filter4[119][2][1] = 35'b00000001001101001101011110110110000;
filter4[119][2][2] = 35'b00001000000111101101011011010000000;
filter4[120][0][0] = 35'b00000001000010100110010000001100000;
filter4[120][0][1] = 35'b11111110001100011010111110100010000;
filter4[120][0][2] = 35'b11111011110010101000100101110000000;
filter4[120][1][0] = 35'b00000100011110000111111000100000000;
filter4[120][1][1] = 35'b11111100010100000111100100100100000;
filter4[120][1][2] = 35'b00000001110101100011110101101000000;
filter4[120][2][0] = 35'b00000011000011101011000101110100000;
filter4[120][2][1] = 35'b00000010010110011011010111111000000;
filter4[120][2][2] = 35'b11111100110000110001100010111000000;
filter4[121][0][0] = 35'b00000010011111010101110000111000000;
filter4[121][0][1] = 35'b11111100111111010000011001101100000;
filter4[121][0][2] = 35'b11111101101101001000010101110100000;
filter4[121][1][0] = 35'b00000011000001001100110101000000000;
filter4[121][1][1] = 35'b00000010000101111111111100000100000;
filter4[121][1][2] = 35'b11111110111101000111011001100010000;
filter4[121][2][0] = 35'b00001001001101100011011101000000000;
filter4[121][2][1] = 35'b00000100011000111110110011111000000;
filter4[121][2][2] = 35'b00000011101110100001110100010000000;
filter4[122][0][0] = 35'b11111111010110101111101000101001000;
filter4[122][0][1] = 35'b11111111111000001001011101011111000;
filter4[122][0][2] = 35'b00000000100010001111001000011101000;
filter4[122][1][0] = 35'b00000000001010010110100001110000010;
filter4[122][1][1] = 35'b00000000010010111101000111001010000;
filter4[122][1][2] = 35'b11111111010001111011110011111000000;
filter4[122][2][0] = 35'b11111101100001110101110101000000000;
filter4[122][2][1] = 35'b11111110000001010001000011110000000;
filter4[122][2][2] = 35'b11110111001111000111000010100000000;
filter4[123][0][0] = 35'b00000000100010010100101111000100000;
filter4[123][0][1] = 35'b11111110101011101111010101000010000;
filter4[123][0][2] = 35'b11111001000000001010100100101000000;
filter4[123][1][0] = 35'b00000010001101110011011010010000000;
filter4[123][1][1] = 35'b00000010100100100011111110110000000;
filter4[123][1][2] = 35'b00000010001100010111010111000000000;
filter4[123][2][0] = 35'b00000010000100111001010100101000000;
filter4[123][2][1] = 35'b00000011000001011111101010101100000;
filter4[123][2][2] = 35'b00000110000100000001011010001000000;
filter4[124][0][0] = 35'b11111111101001010110001101100110100;
filter4[124][0][1] = 35'b00000010101010111100001100001100000;
filter4[124][0][2] = 35'b00000010110001010100111111000100000;
filter4[124][1][0] = 35'b11111100000000100110011101101000000;
filter4[124][1][1] = 35'b11111110001000111000100001010000000;
filter4[124][1][2] = 35'b11111000111100010010010110111000000;
filter4[124][2][0] = 35'b11111110110011011011011101010010000;
filter4[124][2][1] = 35'b11111110011100000011011110101110000;
filter4[124][2][2] = 35'b11111111111111001000000011100010110;
filter4[125][0][0] = 35'b11111001100100110100100111011000000;
filter4[125][0][1] = 35'b11111110011011001000010110001110000;
filter4[125][0][2] = 35'b11111010010111101011011100111000000;
filter4[125][1][0] = 35'b00000001101011001011111001100100000;
filter4[125][1][1] = 35'b00000011011101001010100111110000000;
filter4[125][1][2] = 35'b00000010001001010001111010000000000;
filter4[125][2][0] = 35'b00001000001010010111110111110000000;
filter4[125][2][1] = 35'b00000001000111100000001111100100000;
filter4[125][2][2] = 35'b00000110000100010000011110010000000;
filter4[126][0][0] = 35'b11110110000100010101110000010000000;
filter4[126][0][1] = 35'b11110100101010001100100001100000000;
filter4[126][0][2] = 35'b11111011000110101110100000101000000;
filter4[126][1][0] = 35'b11110001000111011010011011110000000;
filter4[126][1][1] = 35'b11110001011010110010010100010000000;
filter4[126][1][2] = 35'b11111100010000101110000011110000000;
filter4[126][2][0] = 35'b00000000110110100011011001001110000;
filter4[126][2][1] = 35'b11111101101100100010110101001000000;
filter4[126][2][2] = 35'b11111101001101001110111000011100000;
filter4[127][0][0] = 35'b11111100010011111110001111100100000;
filter4[127][0][1] = 35'b11111100001111001111001011111000000;
filter4[127][0][2] = 35'b11111010000011100110000110101000000;
filter4[127][1][0] = 35'b11111011111011011101011100000000000;
filter4[127][1][1] = 35'b11111100010110011100011101010100000;
filter4[127][1][2] = 35'b11111110101011010100011101110000000;
filter4[127][2][0] = 35'b00000011110101101011011000100100000;
filter4[127][2][1] = 35'b00000101100101110110011111101000000;
filter4[127][2][2] = 35'b00000001000011011010011010011000000;

bias4[0] = 35'b00000000001111010011111010011110010;
bias4[1] = 35'b11111110001100001101101000100110000;
bias4[2] = 35'b11111110001110111011001011010100000;
bias4[3] = 35'b11111101011110110011010011010000000;
bias4[4] = 35'b11111100111000100000000110010000000;
bias4[5] = 35'b11111111111000011000000010000010010;
bias4[6] = 35'b00000001100110111111011111011000000;
bias4[7] = 35'b00000010101011101111001101111100000;
bias4[8] = 35'b11111111100111101011001100001110000;
bias4[9] = 35'b00000010010101001111101010000100000;
bias4[10] = 35'b11111101111111010101011010101000000;
bias4[11] = 35'b00000011000100010101000110100100000;
bias4[12] = 35'b00000001001000110011011001000000000;
bias4[13] = 35'b00000011000001110100111000011100000;
bias4[14] = 35'b00000000111001011111111111101010000;
bias4[15] = 35'b00000010111110011001010110110100000;
//================================================================


filter5[0][0] = 35'b00000000011100101110001111001011000;
filter5[0][1] = 35'b00000010111111010010000010000000000;
filter5[0][2] = 35'b11111111110100101000110111100110010;
filter5[0][3] = 35'b11111011110111100011110111000000000;
filter5[0][4] = 35'b11111100110100100011100011110100000;
filter5[0][5] = 35'b00000110101010111000011001101000000;
filter5[0][6] = 35'b00000000001010010100011110111001100;
filter5[0][7] = 35'b11111011100001010101010100001000000;
filter5[0][8] = 35'b11111100011011000101110111011000000;
filter5[0][9] = 35'b00000000110011011010010111101111000;
filter5[0][10] = 35'b00000001000011100011100111100110000;
filter5[0][11] = 35'b00000000010001001010100001100110000;
filter5[0][12] = 35'b00000100100000001011101001111000000;
filter5[0][13] = 35'b11111110001001111001111101000010000;
filter5[0][14] = 35'b00000011001000000011100000111100000;
filter5[0][15] = 35'b00001011011111011101001111000000000;
filter5[0][16] = 35'b11111101100001011111110001111100000;
filter5[0][17] = 35'b11111100000100111011010010100100000;
filter5[0][18] = 35'b00000001001010000011001001000100000;
filter5[0][19] = 35'b11111110010001100100000000010110000;
filter5[0][20] = 35'b00000000100001001001000111000011000;
filter5[0][21] = 35'b11111010000110001101100011000000000;
filter5[0][22] = 35'b00000001111100000011101001111110000;
filter5[0][23] = 35'b00001000000011001001101100000000000;
filter5[0][24] = 35'b00000010100101010101101010001100000;
filter5[0][25] = 35'b11111100011010001101000011001100000;
filter5[0][26] = 35'b11111101101110111110010100010100000;
filter5[0][27] = 35'b11111011100111011101110100001000000;
filter5[0][28] = 35'b11111101011101000001011001110000000;
filter5[0][29] = 35'b11111010010001100000100001001000000;
filter5[0][30] = 35'b00000000011100100010101001001000000;
filter5[0][31] = 35'b00000101000011110111011101100000000;
filter5[0][32] = 35'b00000011101011110001101100110100000;
filter5[0][33] = 35'b11111111111100000000000011000000000;
filter5[0][34] = 35'b00000011000000101101101000101100000;
filter5[0][35] = 35'b00000110001110001111001010001000000;
filter5[0][36] = 35'b11111101000000101000010001111000000;
filter5[0][37] = 35'b00000111010001100000110111011000000;
filter5[0][38] = 35'b11110101100011001001011111110000000;
filter5[0][39] = 35'b00000000001111110011101010111011000;
filter5[0][40] = 35'b11111101011100100111011000001100000;
filter5[0][41] = 35'b00000000010011010100001001101010100;
filter5[0][42] = 35'b11111111110110100001010000110111000;
filter5[0][43] = 35'b11111111111000100011100011000010111;
filter5[0][44] = 35'b00000100110011010000101011000000000;
filter5[0][45] = 35'b00000010110010001110101011011000000;
filter5[0][46] = 35'b11110011011000011011011001010000000;
filter5[0][47] = 35'b11111110010101001000101000100100000;
filter5[0][48] = 35'b00000000010100000010010110011110000;
filter5[0][49] = 35'b11111110000100101101110100010100000;
filter5[0][50] = 35'b11111110101011111100001000011100000;
filter5[0][51] = 35'b00000001101110111110100001100100000;
filter5[0][52] = 35'b00000000111000101000111110101111000;
filter5[0][53] = 35'b00000001101101000100110010011100000;
filter5[0][54] = 35'b11111101011101110110110101000000000;
filter5[0][55] = 35'b11111110110001001111111000000110000;
filter5[0][56] = 35'b00000001001000000110011011001110000;
filter5[0][57] = 35'b11111110110011100100000000001000000;
filter5[0][58] = 35'b11111010100110100111010010000000000;
filter5[0][59] = 35'b00000000001011110011001001010110010;
filter5[0][60] = 35'b11111111100001001010100111010010100;
filter5[0][61] = 35'b11110100011100111110001011010000000;
filter5[0][62] = 35'b11111111010101100010000001111000000;
filter5[0][63] = 35'b00000010110000110001110011000100000;
filter5[0][64] = 35'b11111111000011110101110100011100000;
filter5[0][65] = 35'b11111110110110001100000111011110000;
filter5[0][66] = 35'b00000000011100111101001110101100100;
filter5[0][67] = 35'b11111101101000111010011001100100000;
filter5[0][68] = 35'b11111111100001011011000101101101000;
filter5[0][69] = 35'b00000010011111000000101000000000000;
filter5[0][70] = 35'b00000001010001000110010110011110000;
filter5[0][71] = 35'b11111101101010011111010101111000000;
filter5[0][72] = 35'b11111111000001010001011110000000000;
filter5[0][73] = 35'b11111111111111000101111010000000100;
filter5[0][74] = 35'b00000000001111100001001001011000110;
filter5[0][75] = 35'b11111111101010000011111001010100000;
filter5[0][76] = 35'b00000001011010000000001011101010000;
filter5[0][77] = 35'b00000000010101111011010001110110000;
filter5[0][78] = 35'b11111110000001101010111011000010000;
filter5[0][79] = 35'b00000110001101101011101101000000000;
filter5[0][80] = 35'b11111101000100001000111001100100000;
filter5[0][81] = 35'b11111111001111100111101111011001000;
filter5[0][82] = 35'b11111110111100101101111000111000000;
filter5[0][83] = 35'b00000000100110001011100011011111000;
filter5[0][84] = 35'b11111110111010100100000001010100000;
filter5[0][85] = 35'b11111111110110000001010110100111000;
filter5[0][86] = 35'b11111111100001000011111000111010000;
filter5[0][87] = 35'b00000100011011110110110010110000000;
filter5[0][88] = 35'b11111110010011111010111100100010000;
filter5[0][89] = 35'b11111011001001110110010000011000000;
filter5[0][90] = 35'b11111100110001000101010000110000000;
filter5[0][91] = 35'b11111101101001011011001111011000000;
filter5[0][92] = 35'b11111111010001010001111001010011000;
filter5[0][93] = 35'b11111101010001010001110001100000000;
filter5[0][94] = 35'b11111110000110000110010010010110000;
filter5[0][95] = 35'b00000011001101110110110100010100000;
filter5[0][96] = 35'b00000011100100111010010011010000000;
filter5[0][97] = 35'b11111111111110011111101000000110000;
filter5[0][98] = 35'b00000010000000110011100100110100000;
filter5[0][99] = 35'b00001000010100010111111001000000000;
filter5[0][100] = 35'b11111100010011011000010101011100000;
filter5[0][101] = 35'b00000011010101011001100000010000000;
filter5[0][102] = 35'b11111100010110011101101011001000000;
filter5[0][103] = 35'b11111010000010011101011011011000000;
filter5[0][104] = 35'b11111111111001110110011000110111000;
filter5[0][105] = 35'b11111011011111101111101101111000000;
filter5[0][106] = 35'b00000001110000011110010011010000000;
filter5[0][107] = 35'b00000011110010111001111011001000000;
filter5[0][108] = 35'b00000011100010010001010000110000000;
filter5[0][109] = 35'b11111101110101000101011010001000000;
filter5[0][110] = 35'b00000010001111001010111101101100000;
filter5[0][111] = 35'b11111110011101101100001100100010000;
filter5[0][112] = 35'b00000010110000001001010000000000000;
filter5[0][113] = 35'b11111111010001011100100110010011000;
filter5[0][114] = 35'b11111101000000100100111100001000000;
filter5[0][115] = 35'b11111100011100100101001011101000000;
filter5[0][116] = 35'b11111110101100001001100010110010000;
filter5[0][117] = 35'b00000001001111001000000010110000000;
filter5[0][118] = 35'b00000000110100100011001001111010000;
filter5[0][119] = 35'b00000010011000110000000010010100000;
filter5[0][120] = 35'b11111010011000010011010111100000000;
filter5[0][121] = 35'b00000001000010110100010101110000000;
filter5[0][122] = 35'b00000001010111010000001011001100000;
filter5[0][123] = 35'b11111000110100001111111111000000000;
filter5[0][124] = 35'b11111101110110101011100110010100000;
filter5[0][125] = 35'b11111000011011101101000100101000000;
filter5[0][126] = 35'b11111011100001010001010011111000000;
filter5[0][127] = 35'b00000001010111011100001101011110000;
filter5[0][128] = 35'b11111110101110001111111110100110000;
filter5[0][129] = 35'b11111101101010001011011100000000000;
filter5[0][130] = 35'b11110111010001000001000101010000000;
filter5[0][131] = 35'b11111001110100110001001000011000000;
filter5[0][132] = 35'b00000000101101001100000100100001000;
filter5[0][133] = 35'b00000110010000000100111100111000000;
filter5[0][134] = 35'b00000101000000100010011110101000000;
filter5[0][135] = 35'b11111101100110000100110100000100000;
filter5[0][136] = 35'b11110000110000011110110100100000000;
filter5[0][137] = 35'b11111111110110101011001100000110000;
filter5[0][138] = 35'b11110111110111001111000010010000000;
filter5[0][139] = 35'b11111111110100110101010000101010110;
filter5[0][140] = 35'b00000001101011111011100110101010000;
filter5[0][141] = 35'b11111101100110101110000111000100000;
filter5[0][142] = 35'b11111000101000110110001001110000000;
filter5[0][143] = 35'b00000000010000000000000100111000100;
filter5[0][144] = 35'b11101110111111111111110100100000000;
filter5[0][145] = 35'b11110111110001100000001001000000000;
filter5[0][146] = 35'b11111101011001100011010010001000000;
filter5[0][147] = 35'b00000001000101000010011000101110000;
filter5[0][148] = 35'b00000000101111011010101100110111000;
filter5[0][149] = 35'b00000000010111110001000101011000000;
filter5[0][150] = 35'b00000011011101001100000101111100000;
filter5[0][151] = 35'b11111101100101001110001001110000000;
filter5[0][152] = 35'b11110101111100010001000111010000000;
filter5[0][153] = 35'b11110111011110101110110001100000000;
filter5[0][154] = 35'b00000000011001011000111011000100000;
filter5[0][155] = 35'b11111101111100110101100101101000000;
filter5[0][156] = 35'b00000011011011010111100000011000000;
filter5[0][157] = 35'b11111101011110001110011000001100000;
filter5[0][158] = 35'b11101101011101111110001011100000000;
filter5[0][159] = 35'b11110101010011001000000101010000000;
filter5[0][160] = 35'b11111011010001001010100000111000000;
filter5[0][161] = 35'b11111001110100000101011111111000000;
filter5[0][162] = 35'b00000010010100010111001001101000000;
filter5[0][163] = 35'b00000000011101111000100101110001000;
filter5[0][164] = 35'b00000101011100101100011110101000000;
filter5[0][165] = 35'b11111101100101011100100011001000000;
filter5[0][166] = 35'b11111101100011001000111101110100000;
filter5[0][167] = 35'b11101100011000111000001111100000000;
filter5[0][168] = 35'b11111110000110011111100101100000000;
filter5[0][169] = 35'b00000000010111001100111011010110100;
filter5[0][170] = 35'b11111011101100010001100110011000000;
filter5[0][171] = 35'b00000011011001101100100011001100000;
filter5[0][172] = 35'b00000100110100001110000000100000000;
filter5[0][173] = 35'b11111100000011010100000011110100000;
filter5[0][174] = 35'b00000000101110011101010011101011000;
filter5[0][175] = 35'b11111000101110010010101111010000000;
filter5[0][176] = 35'b00000110101010100000101110000000000;
filter5[0][177] = 35'b11110010100110101011101101000000000;
filter5[0][178] = 35'b11111100011111100110010111001100000;
filter5[0][179] = 35'b00000011111110010010100010110100000;
filter5[0][180] = 35'b00000010000001111101011110111100000;
filter5[0][181] = 35'b11111101001110001110111110111000000;
filter5[0][182] = 35'b11111000100000100100101101101000000;
filter5[0][183] = 35'b11110101111010100001001110000000000;
filter5[0][184] = 35'b11110111101101010101010101010000000;
filter5[0][185] = 35'b11111100011110100001101011001000000;
filter5[0][186] = 35'b11110100011011101100001111010000000;
filter5[0][187] = 35'b11110111100111010000011101010000000;
filter5[0][188] = 35'b11111110101011011101110011100100000;
filter5[0][189] = 35'b11110100111010100101111110110000000;
filter5[0][190] = 35'b11111100111011000100111111111000000;
filter5[0][191] = 35'b11111000011111111111010100101000000;
filter5[0][192] = 35'b00000010110001100101111111000000000;
filter5[0][193] = 35'b11110111001011100010010101110000000;
filter5[0][194] = 35'b00000000111110101111001000110001000;
filter5[0][195] = 35'b11111011111000100111110111101000000;
filter5[0][196] = 35'b11111000111001011011000011100000000;
filter5[0][197] = 35'b11111111110111101000010101101100110;
filter5[0][198] = 35'b11111110100100000100110101111000000;
filter5[0][199] = 35'b11111010000110001100011101111000000;
filter5[0][200] = 35'b11111011101110100010111111110000000;
filter5[0][201] = 35'b11111010100100010110110000000000000;
filter5[0][202] = 35'b11101111110001010100110110100000000;
filter5[0][203] = 35'b00000000011100001101010011011101000;
filter5[0][204] = 35'b11111110000101000011000111101010000;
filter5[0][205] = 35'b00000010000101010111010100000100000;
filter5[0][206] = 35'b00000000001110101011111010100111110;
filter5[0][207] = 35'b11110011011111100010100010100000000;
filter5[0][208] = 35'b11111101101100010000100111011100000;
filter5[0][209] = 35'b11111010000111000010111011110000000;
filter5[0][210] = 35'b11111000110111001011010101000000000;
filter5[0][211] = 35'b11111111110000001010010111010100010;
filter5[0][212] = 35'b00000001001000010000110110011110000;
filter5[0][213] = 35'b00000100000110011000001101011000000;
filter5[0][214] = 35'b11111011001100110110011101110000000;
filter5[0][215] = 35'b11111110001110110101101100011100000;
filter5[0][216] = 35'b11110101110000100000000100010000000;
filter5[0][217] = 35'b11111011100011110000010000100000000;
filter5[0][218] = 35'b00000011010100000011010001111100000;
filter5[0][219] = 35'b11111010000100110110010000000000000;
filter5[0][220] = 35'b11111100010000110000000110001100000;
filter5[0][221] = 35'b11111111000100111110101110010011000;
filter5[0][222] = 35'b00000010110001101100011100110100000;
filter5[0][223] = 35'b00000001100110100001100001010010000;
filter5[0][224] = 35'b11110101111001101111010100000000000;
filter5[0][225] = 35'b11111111010110111010101111001101000;
filter5[0][226] = 35'b11111101100001111011010101011100000;
filter5[0][227] = 35'b00000100110100101100110111000000000;
filter5[0][228] = 35'b00000110010000110000101100110000000;
filter5[0][229] = 35'b11111101110001101010011100110000000;
filter5[0][230] = 35'b11111101010111110001001110111000000;
filter5[0][231] = 35'b11101100010110100011100010000000000;
filter5[0][232] = 35'b11110011001100001111111001010000000;
filter5[0][233] = 35'b11111101000101100011011111000100000;
filter5[0][234] = 35'b11111001011010000100101101010000000;
filter5[0][235] = 35'b00000101011011001011011100010000000;
filter5[0][236] = 35'b11111110111011101001000001000000000;
filter5[0][237] = 35'b11111110011100101000011011001110000;
filter5[0][238] = 35'b11111101011101110111110101000100000;
filter5[0][239] = 35'b11111010000010011001110010100000000;
filter5[0][240] = 35'b11111000001010111111010011100000000;
filter5[0][241] = 35'b00000001000011000000111001010010000;
filter5[0][242] = 35'b11111001101100000001000000010000000;
filter5[0][243] = 35'b00000011100010101100100110111100000;
filter5[0][244] = 35'b00000000001000110111111111001101110;
filter5[0][245] = 35'b00000010100101011000100110110100000;
filter5[0][246] = 35'b11111011110010110011111111000000000;
filter5[0][247] = 35'b00000001000000010001001110000010000;
filter5[0][248] = 35'b11110000001001001111010110010000000;
filter5[0][249] = 35'b00000011000000000111011000111000000;
filter5[0][250] = 35'b11111101110111110111100010011000000;
filter5[0][251] = 35'b00000100011111010011011100101000000;
filter5[0][252] = 35'b11110110100000010110111111010000000;
filter5[0][253] = 35'b00000010010010111101000111001100000;
filter5[0][254] = 35'b11110101010101011100011010100000000;
filter5[0][255] = 35'b11110101001011001001011101010000000;
filter5[0][256] = 35'b00000000110011111110101101101011000;
filter5[0][257] = 35'b11111111001000000001101101011000000;
filter5[0][258] = 35'b11111100011101111110111010110100000;
filter5[0][259] = 35'b11111010010111010000100011100000000;
filter5[0][260] = 35'b11111100110110011101001011001000000;
filter5[0][261] = 35'b11111010010001101011011111111000000;
filter5[0][262] = 35'b11111001011111000100111101111000000;
filter5[0][263] = 35'b11111111000011011100000101001010000;
filter5[0][264] = 35'b11111001001000101011111000100000000;
filter5[0][265] = 35'b11111011101111111101101010001000000;
filter5[0][266] = 35'b11110110011111001101001010110000000;
filter5[0][267] = 35'b11111111111110101100001000001101100;
filter5[0][268] = 35'b11111111111000000010000011110101110;
filter5[0][269] = 35'b00000100001000100001011111000000000;
filter5[0][270] = 35'b11111010100100010011101110010000000;
filter5[0][271] = 35'b11111100000101011011000110001100000;
filter5[0][272] = 35'b11110011011011110011001100100000000;
filter5[0][273] = 35'b11101110100000011001100011000000000;
filter5[0][274] = 35'b11111101100111111011111001111000000;
filter5[0][275] = 35'b00000110100010100101100011100000000;
filter5[0][276] = 35'b00000100110100111000011111011000000;
filter5[0][277] = 35'b11111111100011001001101010011100000;
filter5[0][278] = 35'b11101100000101100100010011000000000;
filter5[0][279] = 35'b11110011101110111011011111100000000;
filter5[0][280] = 35'b11101010011000100100010111000000000;
filter5[0][281] = 35'b11111010101001101001001001111000000;
filter5[0][282] = 35'b11111110001010001101101111100000000;
filter5[0][283] = 35'b00000000001000111000011001011111010;
filter5[0][284] = 35'b00000001001000001001000010111000000;
filter5[0][285] = 35'b11111110001000001001100011010110000;
filter5[0][286] = 35'b00000011010000100111100010001000000;
filter5[0][287] = 35'b11111010010000000010111111001000000;
filter5[0][288] = 35'b00000011111111000101110101011100000;
filter5[0][289] = 35'b11110100010011110000111000010000000;
filter5[0][290] = 35'b11111111001110001101110000100011000;
filter5[0][291] = 35'b11111101111000101110111001110100000;
filter5[0][292] = 35'b00000001100001010001000000100100000;
filter5[0][293] = 35'b11111101111110101000010111110100000;
filter5[0][294] = 35'b11110100111011100011111000110000000;
filter5[0][295] = 35'b11111011100101110110110011110000000;
filter5[0][296] = 35'b11111001000111111110100010101000000;
filter5[0][297] = 35'b00000101010000100101110011100000000;
filter5[0][298] = 35'b00001001111011111011100101100000000;
filter5[0][299] = 35'b11111010110110100010010100100000000;
filter5[0][300] = 35'b00000001011111110100100010111010000;
filter5[0][301] = 35'b11111111111010101110001010001001011;
filter5[0][302] = 35'b00000011001100111000111010011100000;
filter5[0][303] = 35'b11111010100011011110001111110000000;
filter5[0][304] = 35'b11101011100100110110110101000000000;
filter5[0][305] = 35'b00000001111100111101111101100010000;
filter5[0][306] = 35'b11111101100101110111011100010100000;
filter5[0][307] = 35'b11111011111010100000101100100000000;
filter5[0][308] = 35'b00000010000100000010000111100000000;
filter5[0][309] = 35'b00000100110000111101010110011000000;
filter5[0][310] = 35'b11111001011011011010011101110000000;
filter5[0][311] = 35'b11111010010000010011001001111000000;
filter5[0][312] = 35'b11111000100011100111010101010000000;
filter5[0][313] = 35'b11101111100101011001000111100000000;
filter5[0][314] = 35'b00000011110010110101111011000000000;
filter5[0][315] = 35'b11110100110101010001100010110000000;
filter5[0][316] = 35'b00000010110110001101011110111100000;
filter5[0][317] = 35'b11111001001010001000010101001000000;
filter5[0][318] = 35'b11111100101010000011010100010100000;
filter5[0][319] = 35'b11110111011010101111110100100000000;
filter5[0][320] = 35'b00000001110001011010110010001110000;
filter5[0][321] = 35'b00000001100000111101110000010110000;
filter5[0][322] = 35'b00000011000111001000010111110000000;
filter5[0][323] = 35'b00000011111011011001111001111100000;
filter5[0][324] = 35'b00000010100111011010000101011100000;
filter5[0][325] = 35'b00000111011101101111110101000000000;
filter5[0][326] = 35'b00000011001001010101101100010000000;
filter5[0][327] = 35'b00000100100011100001111011011000000;
filter5[0][328] = 35'b11110101111101101000001011010000000;
filter5[0][329] = 35'b11111100001110110101011110010000000;
filter5[0][330] = 35'b11111000100010000000001100011000000;
filter5[0][331] = 35'b00000000010110111101110110101000100;
filter5[0][332] = 35'b00000000010111110010100010011011100;
filter5[0][333] = 35'b11111110110010110100000111011000000;
filter5[0][334] = 35'b00000010011100100001100111001100000;
filter5[0][335] = 35'b00001001100110000100000101110000000;
filter5[0][336] = 35'b11111111001110100101001011110110000;
filter5[0][337] = 35'b11111110001010111101010101010100000;
filter5[0][338] = 35'b11111111011101010111010000000110000;
filter5[0][339] = 35'b11111101101001111000110001100000000;
filter5[0][340] = 35'b00000000011111010111101101111111100;
filter5[0][341] = 35'b00000100110010111011110011011000000;
filter5[0][342] = 35'b00000101111011001011001100110000000;
filter5[0][343] = 35'b00000011000111001010010000111100000;
filter5[0][344] = 35'b00000010011110101110110000011100000;
filter5[0][345] = 35'b11111011101100010011100001111000000;
filter5[0][346] = 35'b00000000001101100110011000010001010;
filter5[0][347] = 35'b11111101110011011010110000011000000;
filter5[0][348] = 35'b11111111000101101000111101110111000;
filter5[0][349] = 35'b11111110100101011011101011101100000;
filter5[0][350] = 35'b00000000100101110100101000100101000;
filter5[0][351] = 35'b00000010011001100101101001110000000;
filter5[0][352] = 35'b11111111000110000011011100110110000;
filter5[0][353] = 35'b00000000001101100010110000011000110;
filter5[0][354] = 35'b00000110011100111001000000111000000;
filter5[0][355] = 35'b11111101011100000101000010110100000;
filter5[0][356] = 35'b11111110110000110101000000001100000;
filter5[0][357] = 35'b00000110010010010011111001101000000;
filter5[0][358] = 35'b11110101100000100111010100000000000;
filter5[0][359] = 35'b11110110101101101110100100110000000;
filter5[0][360] = 35'b00000001011101001100001000001110000;
filter5[0][361] = 35'b11111110000100110110011010111110000;
filter5[0][362] = 35'b11111010000011100001010111000000000;
filter5[0][363] = 35'b00000010010110110100010111101000000;
filter5[0][364] = 35'b00000101001011010100101011110000000;
filter5[0][365] = 35'b00000010011111001001100101110100000;
filter5[0][366] = 35'b11111001100100011101101000111000000;
filter5[0][367] = 35'b00000010000100000111110000100000000;
filter5[0][368] = 35'b00000001001001110110110000001100000;
filter5[0][369] = 35'b11111111001011000111000100001111000;
filter5[0][370] = 35'b00000010100100100001001010111100000;
filter5[0][371] = 35'b00000000101000101111001000100000000;
filter5[0][372] = 35'b11111010011111111101001100111000000;
filter5[0][373] = 35'b00000010001100001010000110001100000;
filter5[0][374] = 35'b11111101100011000000100000100100000;
filter5[0][375] = 35'b11111101101000110100010100111100000;
filter5[0][376] = 35'b11111000110111010110111111111000000;
filter5[0][377] = 35'b11111010111011111111101001111000000;
filter5[0][378] = 35'b11110101011100111100111111000000000;
filter5[0][379] = 35'b11111100110100111000000001110000000;
filter5[0][380] = 35'b11111010110010111010110101110000000;
filter5[0][381] = 35'b11111110101011110100100101111000000;
filter5[0][382] = 35'b00000000101101101110010101100101000;
filter5[0][383] = 35'b11110110011010011010001000110000000;
filter5[0][384] = 35'b11111111010110001011010001110000000;
filter5[0][385] = 35'b11111111111001111010001010001111001;
filter5[0][386] = 35'b00000000101011010001101000011000000;
filter5[0][387] = 35'b11111110101011000100101000011110000;
filter5[0][388] = 35'b11111110111101000111000001101100000;
filter5[0][389] = 35'b11111110101101100011111101001000000;
filter5[0][390] = 35'b11111111100010001101111110010001100;
filter5[0][391] = 35'b00000001111110111011110111001100000;
filter5[0][392] = 35'b11111110110011000010101111001110000;
filter5[0][393] = 35'b00000000011011111001010000110001000;
filter5[0][394] = 35'b11111110110010111000000000110000000;
filter5[0][395] = 35'b00000000100110111101101101001010000;
filter5[0][396] = 35'b00000000010011111010101001101001000;
filter5[0][397] = 35'b11111111011000100010111010001011000;
filter5[0][398] = 35'b00000010000100001001001010110100000;
filter5[0][399] = 35'b00000011000110101000000001101100000;
filter5[0][400] = 35'b11111111101111001111011010001100000;
filter5[0][401] = 35'b00000000011011010110110110001101000;
filter5[0][402] = 35'b11111110111001011011111110010010000;
filter5[0][403] = 35'b11111100111011011100010100001100000;
filter5[0][404] = 35'b00000000001100110101100010101000110;
filter5[0][405] = 35'b00000000110001110001101100001000000;
filter5[0][406] = 35'b00000001110110000000010110011100000;
filter5[0][407] = 35'b00000011000100000001110000001100000;
filter5[0][408] = 35'b00000001010010000011010111000010000;
filter5[0][409] = 35'b00000000011010100010100101010001100;
filter5[0][410] = 35'b00000010010010100100001001101000000;
filter5[0][411] = 35'b00000000101111001100100010111000000;
filter5[0][412] = 35'b11111111010110110011100011010101000;
filter5[0][413] = 35'b11111110110011110100011011100100000;
filter5[0][414] = 35'b11111101100111100110011000000100000;
filter5[0][415] = 35'b00000000100000010010001101011100000;
filter5[0][416] = 35'b11111110001010000001011110100010000;
filter5[0][417] = 35'b11111111101011110000100000011111000;
filter5[0][418] = 35'b00000111100001110100110100010000000;
filter5[0][419] = 35'b00000010110011111111011110010100000;
filter5[0][420] = 35'b00000000010000101111011000111010000;
filter5[0][421] = 35'b11111110000001110000011001000000000;
filter5[0][422] = 35'b00000010000110101010000110101100000;
filter5[0][423] = 35'b11111000010111110101100010111000000;
filter5[0][424] = 35'b11111101001010010101011000100000000;
filter5[0][425] = 35'b00000010110000010011101001111000000;
filter5[0][426] = 35'b11111100100101000010001100111100000;
filter5[0][427] = 35'b11111101110000101100001110011000000;
filter5[0][428] = 35'b00000111111010000101111011110000000;
filter5[0][429] = 35'b00000001010100011011100010101010000;
filter5[0][430] = 35'b00000010100001010101100100111100000;
filter5[0][431] = 35'b11111110011101111111001100101010000;
filter5[0][432] = 35'b11111111000010100100101001100111000;
filter5[0][433] = 35'b11111011001110010001100001001000000;
filter5[0][434] = 35'b11111111001101010101111010101101000;
filter5[0][435] = 35'b11111101011010111101000001100000000;
filter5[0][436] = 35'b11111100000101110011101110101100000;
filter5[0][437] = 35'b00000110011100000111000110011000000;
filter5[0][438] = 35'b11111011111100001101101100010000000;
filter5[0][439] = 35'b00000000001100100100001111110110110;
filter5[0][440] = 35'b11111101001110010001011010111100000;
filter5[0][441] = 35'b11111111110011110000101011111101010;
filter5[0][442] = 35'b00000001011001001010011100101010000;
filter5[0][443] = 35'b00000000011001001011100000011111100;
filter5[0][444] = 35'b11111101000101010111001100000100000;
filter5[0][445] = 35'b11111111111010001111100111011111101;
filter5[0][446] = 35'b00000000111011111001000111101101000;
filter5[0][447] = 35'b00000000111110101110111011101011000;
filter5[0][448] = 35'b00000001000011110111010010100000000;
filter5[0][449] = 35'b11111111001101010001101100100100000;
filter5[0][450] = 35'b11111011010110111000110101101000000;
filter5[0][451] = 35'b00000011010101001110111101011000000;
filter5[0][452] = 35'b00000000110011101101001110000001000;
filter5[0][453] = 35'b11111111011011010001001001101101000;
filter5[0][454] = 35'b00000000001000011011010111000111110;
filter5[0][455] = 35'b11111100100001001101011101000100000;
filter5[0][456] = 35'b11111111100001101101111100100010100;
filter5[0][457] = 35'b00000001001111000111001100010110000;
filter5[0][458] = 35'b11111111111111011011101000110111001;
filter5[0][459] = 35'b00000011101011000000111000110000000;
filter5[0][460] = 35'b00000010111011100010001010010000000;
filter5[0][461] = 35'b00000011101011001001101110000100000;
filter5[0][462] = 35'b00000110111111000100101010100000000;
filter5[0][463] = 35'b11111101010000001100011110001100000;
filter5[0][464] = 35'b11111011011010100000100101100000000;
filter5[0][465] = 35'b00000101111110011111011011111000000;
filter5[0][466] = 35'b11111101011110010011101110110100000;
filter5[0][467] = 35'b11111000010110110111100110111000000;
filter5[0][468] = 35'b11111110101001101100101101010010000;
filter5[0][469] = 35'b00001010011111100011110100010000000;
filter5[0][470] = 35'b11111110110010100010011110100100000;
filter5[0][471] = 35'b00000101101110000110011111011000000;
filter5[0][472] = 35'b11110111100101101010010000010000000;
filter5[0][473] = 35'b00000001110001110010001011110010000;
filter5[0][474] = 35'b00000001000010101001010011101000000;
filter5[0][475] = 35'b11111111100111110111101101000110000;
filter5[0][476] = 35'b11111101010101101110100000101000000;
filter5[0][477] = 35'b11111101000001001000110000101100000;
filter5[0][478] = 35'b11111111011010011100101100111010000;
filter5[0][479] = 35'b00000100011011100110000100011000000;
filter5[0][480] = 35'b11111010111011011010100101101000000;
filter5[0][481] = 35'b00000001100011100000100111011000000;
filter5[0][482] = 35'b00000010110010111110011001110000000;
filter5[0][483] = 35'b11111110011111001010100111110010000;
filter5[0][484] = 35'b00000101101000110100010111111000000;
filter5[0][485] = 35'b00000000011001110110010000110001000;
filter5[0][486] = 35'b11111101111110011101001000110000000;
filter5[0][487] = 35'b11111001111011110111111000000000000;
filter5[0][488] = 35'b00001000000111001011000010010000000;
filter5[0][489] = 35'b11111101100010010111010100110100000;
filter5[0][490] = 35'b00000001100010111100110101000110000;
filter5[0][491] = 35'b11111111011010010000110000100010000;
filter5[0][492] = 35'b00000000001000101010010011111011100;
filter5[0][493] = 35'b11111110000111100011011111111100000;
filter5[0][494] = 35'b11111101101011100010001001001100000;
filter5[0][495] = 35'b11110011000011110001110000110000000;
filter5[0][496] = 35'b00000011101101010000010001000100000;
filter5[0][497] = 35'b11111011100110110110100001000000000;
filter5[0][498] = 35'b11111111011101000110101010100011000;
filter5[0][499] = 35'b00000000100111110011100110000000000;
filter5[0][500] = 35'b00000100000000011011011101100000000;
filter5[0][501] = 35'b00000001001001010101011010101000000;
filter5[0][502] = 35'b11111110100010100000100100100000000;
filter5[0][503] = 35'b00000000111110011010100010100010000;
filter5[0][504] = 35'b11111011000111111101010010011000000;
filter5[0][505] = 35'b11111111111110111101010010100000011;
filter5[0][506] = 35'b00000000010100110101111101000100100;
filter5[0][507] = 35'b00000000010010111111001001001011000;
filter5[0][508] = 35'b11111101110011100101010011100000000;
filter5[0][509] = 35'b00000100010001101110000001101000000;
filter5[0][510] = 35'b11111101110010001111110000010000000;
filter5[0][511] = 35'b00000000000100000111110101001110110;
filter5[0][512] = 35'b11111110001110100001111111001010000;
filter5[0][513] = 35'b11111111000110101101011101001010000;
filter5[0][514] = 35'b11111111111001000110100100011110010;
filter5[0][515] = 35'b11111100110101101010000100001000000;
filter5[0][516] = 35'b00000011010011101110011011010100000;
filter5[0][517] = 35'b00000011000011000010101101111000000;
filter5[0][518] = 35'b00000100110001011101000010011000000;
filter5[0][519] = 35'b00000100001010000010011010010000000;
filter5[0][520] = 35'b11111111110010000001110111110111000;
filter5[0][521] = 35'b11111100111111011101111101100000000;
filter5[0][522] = 35'b11111011111100011000000111111000000;
filter5[0][523] = 35'b11111101111111100110011101010000000;
filter5[0][524] = 35'b00000001000001011001101001100010000;
filter5[0][525] = 35'b11111111000001000100100010000100000;
filter5[0][526] = 35'b11111110111010101001110111100100000;
filter5[0][527] = 35'b00000110001101001100011010110000000;
filter5[0][528] = 35'b11111101110011000011110101011100000;
filter5[0][529] = 35'b00000000110001110101100010100011000;
filter5[0][530] = 35'b11111111101000000110000101011111100;
filter5[0][531] = 35'b11111010010011101111100001011000000;
filter5[0][532] = 35'b11111111010001000110111001101000000;
filter5[0][533] = 35'b00000110000110111101110110010000000;
filter5[0][534] = 35'b11111111000010111000110111010101000;
filter5[0][535] = 35'b00000010011110101111101100001100000;
filter5[0][536] = 35'b11111101000000110000010100001000000;
filter5[0][537] = 35'b11111110010011001001100000111000000;
filter5[0][538] = 35'b11111111100101000110100011100010000;
filter5[0][539] = 35'b00000100001001101010111001110000000;
filter5[0][540] = 35'b11111110001111100100010111000110000;
filter5[0][541] = 35'b00000010001111010110000011000000000;
filter5[0][542] = 35'b11111111110011010001101100000111100;
filter5[0][543] = 35'b00000000011110001000001110101010100;
filter5[0][544] = 35'b00000000011001111110110101011110100;
filter5[0][545] = 35'b00000000111111010010001101010001000;
filter5[0][546] = 35'b00000100010110110010000100110000000;
filter5[0][547] = 35'b11111101000000000101000011011100000;
filter5[0][548] = 35'b11111101001111011111100101000000000;
filter5[0][549] = 35'b00000001011100100110100100100110000;
filter5[0][550] = 35'b11111100011100110100010110101100000;
filter5[0][551] = 35'b11111111100010011011111110100101000;
filter5[0][552] = 35'b00000000010011001001001011110111100;
filter5[0][553] = 35'b00000001101111010101110110001010000;
filter5[0][554] = 35'b11111010111011011101100111011000000;
filter5[0][555] = 35'b00000000110100001011010101001011000;
filter5[0][556] = 35'b00000111100001101100101001000000000;
filter5[0][557] = 35'b00000010010001011101011110100000000;
filter5[0][558] = 35'b11111100001111110010011100001100000;
filter5[0][559] = 35'b11111100100001001000101001110100000;
filter5[0][560] = 35'b11111110001110110011111010101100000;
filter5[0][561] = 35'b00000001100010001101100000011110000;
filter5[0][562] = 35'b11111101101010111110001001010100000;
filter5[0][563] = 35'b00000000111100111110110111011011000;
filter5[0][564] = 35'b11111101111110110110101010100000000;
filter5[0][565] = 35'b00000001100110010011111100111000000;
filter5[0][566] = 35'b00000101111110101001010100111000000;
filter5[0][567] = 35'b11111111000001010110010100101000000;
filter5[0][568] = 35'b11111110101011000001110000001000000;
filter5[0][569] = 35'b11111100010011100011111010101000000;
filter5[0][570] = 35'b00000011001100001010100110000100000;
filter5[0][571] = 35'b11111111000000010101001011001001000;
filter5[0][572] = 35'b11111101110001110101010110011000000;
filter5[0][573] = 35'b11111101000101111101010100010000000;
filter5[0][574] = 35'b00000000010011000101110110010010100;
filter5[0][575] = 35'b00000011000000010011010000000100000;
filter5[0][576] = 35'b11111111010101110010110010111010000;
filter5[0][577] = 35'b00000010111011001010010100110000000;
filter5[0][578] = 35'b11111100111111110110101011000100000;
filter5[0][579] = 35'b00000000111011000011100110010000000;
filter5[0][580] = 35'b11111111001101001101111001010001000;
filter5[0][581] = 35'b00000010101010111101011100100100000;
filter5[0][582] = 35'b00000100111000100110111001110000000;
filter5[0][583] = 35'b00000100000000000100011110100000000;
filter5[0][584] = 35'b00000000001001110111001100110111110;
filter5[0][585] = 35'b11111110000101011111000000100110000;
filter5[0][586] = 35'b11111100100100001111000111000100000;
filter5[0][587] = 35'b11111011001100001011101100111000000;
filter5[0][588] = 35'b11111111101100001111000101000111100;
filter5[0][589] = 35'b11111111100000101100010110011110000;
filter5[0][590] = 35'b00000001100011010000011000010000000;
filter5[0][591] = 35'b11111110010011000010000010110110000;
filter5[0][592] = 35'b11111101011100000011001010010100000;
filter5[0][593] = 35'b00000010011110000001110001010100000;
filter5[0][594] = 35'b11111101000011111000010000101100000;
filter5[0][595] = 35'b11111101110101101010101101001100000;
filter5[0][596] = 35'b11111101000101100110000111100000000;
filter5[0][597] = 35'b00000000110110000011100100100111000;
filter5[0][598] = 35'b11111111101000010000100010011000100;
filter5[0][599] = 35'b00000000000110100101100111111110011;
filter5[0][600] = 35'b11111010011000001101001001001000000;
filter5[0][601] = 35'b00000000000011101001000101010011110;
filter5[0][602] = 35'b11111111100001110010010001101110100;
filter5[0][603] = 35'b00000100001100100111010100011000000;
filter5[0][604] = 35'b11111110111010011001110100011110000;
filter5[0][605] = 35'b00000001010110100110100011011000000;
filter5[0][606] = 35'b11111101100110011001111010111100000;
filter5[0][607] = 35'b11111100111111011100101110111000000;
filter5[0][608] = 35'b11111110100000110111000010011100000;
filter5[0][609] = 35'b11111111011011001011010010010100000;
filter5[0][610] = 35'b00000001111001111101111011010000000;
filter5[0][611] = 35'b00000101001001010001100011000000000;
filter5[0][612] = 35'b00000010000011101101000110010100000;
filter5[0][613] = 35'b11111110100001110111110000111000000;
filter5[0][614] = 35'b11111101111001110011011011000100000;
filter5[0][615] = 35'b11111011010101000110011001100000000;
filter5[0][616] = 35'b11111110001111010010110010111000000;
filter5[0][617] = 35'b00000100000101011010101010100000000;
filter5[0][618] = 35'b11110111000011000111110000100000000;
filter5[0][619] = 35'b11111111011100111001110000010000000;
filter5[0][620] = 35'b00000101110001001011001110111000000;
filter5[0][621] = 35'b00000010110111100011011011111100000;
filter5[0][622] = 35'b11111110000001010000010111111010000;
filter5[0][623] = 35'b00000010111111101010001111101100000;
filter5[0][624] = 35'b11111101101011000110001000110100000;
filter5[0][625] = 35'b11111010001101000011101011000000000;
filter5[0][626] = 35'b11111000000001101100000110000000000;
filter5[0][627] = 35'b11111110100000001001011011010110000;
filter5[0][628] = 35'b00000000111001100101100000111011000;
filter5[0][629] = 35'b00000100110111110010000101100000000;
filter5[0][630] = 35'b00000001101111001011010101011100000;
filter5[0][631] = 35'b11111111111110000111001000110000101;
filter5[0][632] = 35'b00000001010010011010000001011010000;
filter5[0][633] = 35'b00001001100001011011111001000000000;
filter5[0][634] = 35'b00000010001001000111001101001100000;
filter5[0][635] = 35'b11111100100011101101010000010100000;
filter5[0][636] = 35'b11111010000000111100001100011000000;
filter5[0][637] = 35'b11111101110011000011010101000000000;
filter5[0][638] = 35'b11111000100101001110011011100000000;
filter5[0][639] = 35'b11111111010101100110000011001111000;
filter5[0][640] = 35'b00000001110100110000101100001010000;
filter5[0][641] = 35'b11111101001010101001110011010000000;
filter5[0][642] = 35'b00000001011100000101010101101000000;
filter5[0][643] = 35'b11111110101000010001100101000110000;
filter5[0][644] = 35'b11111100001000101000101110101000000;
filter5[0][645] = 35'b00000010110100000000101011110100000;
filter5[0][646] = 35'b00000000101010111000000110001001000;
filter5[0][647] = 35'b11111100110000111111010110000100000;
filter5[0][648] = 35'b00000001011010100011101000010110000;
filter5[0][649] = 35'b00000010110110011010101101100100000;
filter5[0][650] = 35'b00000010001001010111100001001000000;
filter5[0][651] = 35'b11111101100001111001100000000100000;
filter5[0][652] = 35'b00000000111010110011011101010011000;
filter5[0][653] = 35'b00000001110011010010110010111000000;
filter5[0][654] = 35'b00000010011001111010100101110100000;
filter5[0][655] = 35'b00000101001111000101101110101000000;
filter5[0][656] = 35'b11111100011111010110011000001100000;
filter5[0][657] = 35'b11111110101101011000101110001110000;
filter5[0][658] = 35'b11111100110011110100110110111100000;
filter5[0][659] = 35'b11111000111110001010010110101000000;
filter5[0][660] = 35'b11111100100010101101111110101000000;
filter5[0][661] = 35'b00000001100100011010011001101110000;
filter5[0][662] = 35'b00000000000101100001000000110101100;
filter5[0][663] = 35'b00000101100101001111001000100000000;
filter5[0][664] = 35'b00000010111000111010000110001000000;
filter5[0][665] = 35'b11111010111001000100001011110000000;
filter5[0][666] = 35'b11111101110111111010101101001100000;
filter5[0][667] = 35'b11111111011101010101011000010011000;
filter5[0][668] = 35'b11111010100110101101000000000000000;
filter5[0][669] = 35'b11111100001111011100101110101000000;
filter5[0][670] = 35'b11111011101110110110101111010000000;
filter5[0][671] = 35'b00000100010111001111100100000000000;
filter5[0][672] = 35'b00000010111111010111110111100100000;
filter5[0][673] = 35'b00000001011111001000001010011110000;
filter5[0][674] = 35'b11111011111110111010100111010000000;
filter5[0][675] = 35'b11111101000101010011001111000000000;
filter5[0][676] = 35'b00000100001001111111101100110000000;
filter5[0][677] = 35'b11111111001110100010010000110101000;
filter5[0][678] = 35'b11111111101111110101010011110110000;
filter5[0][679] = 35'b11111101011110011101110000000000000;
filter5[0][680] = 35'b11111101111001110101111000100100000;
filter5[0][681] = 35'b00000100111000010101011110111000000;
filter5[0][682] = 35'b00000001111110000000010010000010000;
filter5[0][683] = 35'b11111111010011111101110010011001000;
filter5[0][684] = 35'b00000010001110111110010110111000000;
filter5[0][685] = 35'b00000010111110010010011101010000000;
filter5[0][686] = 35'b00000000000011110111111101000100100;
filter5[0][687] = 35'b11110111000011001101000110110000000;
filter5[0][688] = 35'b00000001011101110011010011010000000;
filter5[0][689] = 35'b00000001111010011001011110011110000;
filter5[0][690] = 35'b11111000101001100101100011010000000;
filter5[0][691] = 35'b00000011100000110000010000011000000;
filter5[0][692] = 35'b00000101110100111110100011110000000;
filter5[0][693] = 35'b11111100110111111111101100011100000;
filter5[0][694] = 35'b00000011000001011011110110100100000;
filter5[0][695] = 35'b11111111000010000011010001000110000;
filter5[0][696] = 35'b11111101101011111100010110111100000;
filter5[0][697] = 35'b11111101101100001101000101000000000;
filter5[0][698] = 35'b11111100011101001100011001000100000;
filter5[0][699] = 35'b00000001000111110100001100111000000;
filter5[0][700] = 35'b11111110100101100100001001111010000;
filter5[0][701] = 35'b00000001111001001010111110001010000;
filter5[0][702] = 35'b11111111101110010010100001010011000;
filter5[0][703] = 35'b00000001111111100000001110010100000;
filter5[0][704] = 35'b00000000010111010100101110111011100;
filter5[0][705] = 35'b11111111011110011101010000000100000;
filter5[0][706] = 35'b11111111001011101010010011101110000;
filter5[0][707] = 35'b11111110011111010010111011101010000;
filter5[0][708] = 35'b11111111111011101111111001010101111;
filter5[0][709] = 35'b00000000100001001111001001100001000;
filter5[0][710] = 35'b11111110110111000100111010110100000;
filter5[0][711] = 35'b11111111010110100000010010100001000;
filter5[0][712] = 35'b11111110011010101110101011110100000;
filter5[0][713] = 35'b00000001000010011100001010111100000;
filter5[0][714] = 35'b11111111110100001011111100010110110;
filter5[0][715] = 35'b00000001000001011011010010010000000;
filter5[0][716] = 35'b11111111110011011111100001101000000;
filter5[0][717] = 35'b00000001011010001100100100110110000;
filter5[0][718] = 35'b00000000100111010110010001100000000;
filter5[0][719] = 35'b11111111000101010100111110010011000;
filter5[0][720] = 35'b00000000111001101100110110111001000;
filter5[0][721] = 35'b11111111101111110110111001100011000;
filter5[0][722] = 35'b11111111101000010101110000010010100;
filter5[0][723] = 35'b00000001010011001010111110000010000;
filter5[0][724] = 35'b00000001011110100100010101110100000;
filter5[0][725] = 35'b00000001000010000000011110101000000;
filter5[0][726] = 35'b00000001100100110010011000100000000;
filter5[0][727] = 35'b00000000100111011100100011100000000;
filter5[0][728] = 35'b11111110110110111110110011110000000;
filter5[0][729] = 35'b11111110010111010100100110000000000;
filter5[0][730] = 35'b00000000001101111000001101110011100;
filter5[0][731] = 35'b11111101000100110100101101101000000;
filter5[0][732] = 35'b00000000101000011001000101110011000;
filter5[0][733] = 35'b11111110001100011101101111110000000;
filter5[0][734] = 35'b00000000110111100010000101000111000;
filter5[0][735] = 35'b11111110011100101010000101011000000;
filter5[0][736] = 35'b11111111010101001110000100011001000;
filter5[0][737] = 35'b11111010111010101011000111001000000;
filter5[0][738] = 35'b00000000111010101110001100000100000;
filter5[0][739] = 35'b11111111010011010011010101000011000;
filter5[0][740] = 35'b00000000101110010111101100111000000;
filter5[0][741] = 35'b11111101101101000000011000010100000;
filter5[0][742] = 35'b11111101011100011110101110000000000;
filter5[0][743] = 35'b11111110010101001111110001010110000;
filter5[0][744] = 35'b11111101110011100101101011000000000;
filter5[0][745] = 35'b11111010011100001100111001100000000;
filter5[0][746] = 35'b11111101110010101001101101001100000;
filter5[0][747] = 35'b00000011001111111001110010001000000;
filter5[0][748] = 35'b00000101000100100000010110010000000;
filter5[0][749] = 35'b00000010101110110101101011000100000;
filter5[0][750] = 35'b11111100111011011111000110011100000;
filter5[0][751] = 35'b00000010110011001100110001000000000;
filter5[0][752] = 35'b11111101110111111111001100000100000;
filter5[0][753] = 35'b00000011000100010011100100100000000;
filter5[0][754] = 35'b11111001011111111110101100000000000;
filter5[0][755] = 35'b00000100000100010011011110110000000;
filter5[0][756] = 35'b00000010101010101100001101011100000;
filter5[0][757] = 35'b11111101110100011111101011010100000;
filter5[0][758] = 35'b11111100001100110110000001001000000;
filter5[0][759] = 35'b11111110001101110011100100111110000;
filter5[0][760] = 35'b11111110110011101010000100101010000;
filter5[0][761] = 35'b00000000110001111001010101010111000;
filter5[0][762] = 35'b00000000000001011000010111001000110;
filter5[0][763] = 35'b00000001111101011011111111100010000;
filter5[0][764] = 35'b11111100001110100010100110111000000;
filter5[0][765] = 35'b11111110101110101001010001010100000;
filter5[0][766] = 35'b00000000011101101010101100001000000;
filter5[0][767] = 35'b11111101101101000100000110001100000;
filter5[0][768] = 35'b11111100100010100100001001011000000;
filter5[0][769] = 35'b11111110111101001110011100110010000;
filter5[0][770] = 35'b11111110110000010000010011111100000;
filter5[0][771] = 35'b11111110000011111011010001111110000;
filter5[0][772] = 35'b00000001101011001100011100100100000;
filter5[0][773] = 35'b11111111111010011100111111011000000;
filter5[0][774] = 35'b00000001100011000100001101011000000;
filter5[0][775] = 35'b00000011011000111110101100011000000;
filter5[0][776] = 35'b11111101010100000111010011011100000;
filter5[0][777] = 35'b11111111100001000001010100100000000;
filter5[0][778] = 35'b11111111110001111101001001111001110;
filter5[0][779] = 35'b11111110111111100000001011010010000;
filter5[0][780] = 35'b00000000000011000111001001111010010;
filter5[0][781] = 35'b00000010010001001101101001010000000;
filter5[0][782] = 35'b00000010110010111010010010110100000;
filter5[0][783] = 35'b11111100000111111011011001101100000;
filter5[0][784] = 35'b11111110111111101000001101010000000;
filter5[0][785] = 35'b11111110101001000100000110011100000;
filter5[0][786] = 35'b11111111011110101010011100110010000;
filter5[0][787] = 35'b11111110000001101100110111001000000;
filter5[0][788] = 35'b00000001001100110001011010001010000;
filter5[0][789] = 35'b00000001110011010100000110001110000;
filter5[0][790] = 35'b00000000100101111011001010011110000;
filter5[0][791] = 35'b11111111000011111110000011110010000;
filter5[0][792] = 35'b11111001010001011100010100110000000;
filter5[0][793] = 35'b00000000101010010011100010010000000;
filter5[0][794] = 35'b11111011110111101111111111001000000;
filter5[0][795] = 35'b11111111101101010000110110100101000;
filter5[0][796] = 35'b11111111010011000010001111011011000;
filter5[0][797] = 35'b00000100111110100010010110111000000;
filter5[0][798] = 35'b11111000111100101000100111111000000;
filter5[0][799] = 35'b00000010100100010110111011100000000;
filter5[0][800] = 35'b11111111100110010001101010100110000;
filter5[0][801] = 35'b11111111011100011111001001101110000;
filter5[0][802] = 35'b00000010111111110101010011001100000;
filter5[0][803] = 35'b00000010100110001101100111000000000;
filter5[0][804] = 35'b11111110101001111100110000100010000;
filter5[0][805] = 35'b11111111011110010100011101000001000;
filter5[0][806] = 35'b11111110101001011001101101100110000;
filter5[0][807] = 35'b11111101001000000100001010000000000;
filter5[0][808] = 35'b00000000001011010101000111001111010;
filter5[0][809] = 35'b11111001010011001010010001110000000;
filter5[0][810] = 35'b11111011100011011101101010001000000;
filter5[0][811] = 35'b00000101100101111001100100110000000;
filter5[0][812] = 35'b11111110000011010000000010101100000;
filter5[0][813] = 35'b00000010111000111100110110011000000;
filter5[0][814] = 35'b00000001001011111000100001011100000;
filter5[0][815] = 35'b11111110101001101011001000000000000;
filter5[0][816] = 35'b00000001101100011101000100111110000;
filter5[0][817] = 35'b11111111001011010000010011110111000;
filter5[0][818] = 35'b11111111110010111101011001010101110;
filter5[0][819] = 35'b00001000010000110101100111010000000;
filter5[0][820] = 35'b00000011101000111101010011000100000;
filter5[0][821] = 35'b11111111011101110100101101011111000;
filter5[0][822] = 35'b11111100100100101100011000000000000;
filter5[0][823] = 35'b11111101111101100000001011110100000;
filter5[0][824] = 35'b00000001101100111101011110011010000;
filter5[0][825] = 35'b11111101001001001011101100110000000;
filter5[0][826] = 35'b11110111100101000111110110010000000;
filter5[0][827] = 35'b00000111001100100100001100110000000;
filter5[0][828] = 35'b11111111010111001010001111101101000;
filter5[0][829] = 35'b00000010101110011010011110110000000;
filter5[0][830] = 35'b00000010010000101100000100110100000;
filter5[0][831] = 35'b11111111011111001111000001001001000;
filter5[0][832] = 35'b11111110011111111111011110111100000;
filter5[0][833] = 35'b00000000100000111011000000101110000;
filter5[0][834] = 35'b11111111011011111010111110001100000;
filter5[0][835] = 35'b11111111110010111001001011011010000;
filter5[0][836] = 35'b11111111101001100101110111011001100;
filter5[0][837] = 35'b11111110101001110111001110010010000;
filter5[0][838] = 35'b11111111111111010100001000001101000;
filter5[0][839] = 35'b11111111001111110110011001010110000;
filter5[0][840] = 35'b00000000100100111000110101100111000;
filter5[0][841] = 35'b11111111100111100000000011100100000;
filter5[0][842] = 35'b11111111111001111100000100100010100;
filter5[0][843] = 35'b11111110111110101111010001100110000;
filter5[0][844] = 35'b11111111001100111010110010111000000;
filter5[0][845] = 35'b11111111111000010100101111101101101;
filter5[0][846] = 35'b11111111101000000010010011001011100;
filter5[0][847] = 35'b00000000110010100011011101010100000;
filter5[0][848] = 35'b11111111001110011100110001110000000;
filter5[0][849] = 35'b11111110111011011010001111000110000;
filter5[0][850] = 35'b11111111001000110101010110001100000;
filter5[0][851] = 35'b11111111100111111110111101001110000;
filter5[0][852] = 35'b00000000111011111010111011001110000;
filter5[0][853] = 35'b00000000001110000011000100001000100;
filter5[0][854] = 35'b11111101110000100111001111000000000;
filter5[0][855] = 35'b11111111011001101000000100011000000;
filter5[0][856] = 35'b11111111011101001110001100100010000;
filter5[0][857] = 35'b00000000001001011001010100100001010;
filter5[0][858] = 35'b11111101111010110011000110011100000;
filter5[0][859] = 35'b00000000100001110110100110110000000;
filter5[0][860] = 35'b11111110010100010111001011100110000;
filter5[0][861] = 35'b11111101111100110101000111000100000;
filter5[0][862] = 35'b00000010110011110111011110110100000;
filter5[0][863] = 35'b00000000011101110100000010001000000;
filter5[0][864] = 35'b11111110100000000100100110110100000;
filter5[0][865] = 35'b00000000000011100001011001010111001;
filter5[0][866] = 35'b11111100101100000010100000110100000;
filter5[0][867] = 35'b00000001010111010010011011001010000;
filter5[0][868] = 35'b00000000100111011000101101101011000;
filter5[0][869] = 35'b11111110110101100000000001101010000;
filter5[0][870] = 35'b11111011110110000100101101101000000;
filter5[0][871] = 35'b00000010000000111010000011100100000;
filter5[0][872] = 35'b00000000000110101011111000001100001;
filter5[0][873] = 35'b11111100110011110000110010110100000;
filter5[0][874] = 35'b00000010100001001001010011001000000;
filter5[0][875] = 35'b00000100111001010011110111110000000;
filter5[0][876] = 35'b11111010010101000001000001000000000;
filter5[0][877] = 35'b11111100111111110001111110111100000;
filter5[0][878] = 35'b11111110101100110011001010000000000;
filter5[0][879] = 35'b11111101011111011011000111111100000;
filter5[0][880] = 35'b00000000010111101111000000101010000;
filter5[0][881] = 35'b00000000001000110100101010110010100;
filter5[0][882] = 35'b11111101111010100111101100110100000;
filter5[0][883] = 35'b00000101011000100011000100001000000;
filter5[0][884] = 35'b00000101110101100010000100000000000;
filter5[0][885] = 35'b11111100001100000110010100000000000;
filter5[0][886] = 35'b00000100000111010100100111011000000;
filter5[0][887] = 35'b11111111001111000101001010000000000;
filter5[0][888] = 35'b11111101010100100001001001001100000;
filter5[0][889] = 35'b11111101110010001101101101011100000;
filter5[0][890] = 35'b00000000110000111100011011011111000;
filter5[0][891] = 35'b11111100100010101001000100110000000;
filter5[0][892] = 35'b11111111100110000011110011011101100;
filter5[0][893] = 35'b00000001001001011001010010111000000;
filter5[0][894] = 35'b00000010010111010010110010100000000;
filter5[0][895] = 35'b00000000111100110001110100111101000;
filter5[0][896] = 35'b11111101110100100010100111111000000;
filter5[0][897] = 35'b00000001110011101110111111000100000;
filter5[0][898] = 35'b00000010101011101110111101001100000;
filter5[0][899] = 35'b11110001110101111111000100010000000;
filter5[0][900] = 35'b00000001001100001111110001100010000;
filter5[0][901] = 35'b00001000010011110011010101100000000;
filter5[0][902] = 35'b11110110111010011000001101100000000;
filter5[0][903] = 35'b11111011101111011000010110000000000;
filter5[0][904] = 35'b11111001111100001011001110010000000;
filter5[0][905] = 35'b11111101100001000100111110110000000;
filter5[0][906] = 35'b11111001101101110000011110011000000;
filter5[0][907] = 35'b11111010001011001010111000000000000;
filter5[0][908] = 35'b11111111100010011111100110101100100;
filter5[0][909] = 35'b00000100101100101100100010111000000;
filter5[0][910] = 35'b11110110101011011110100000110000000;
filter5[0][911] = 35'b11111100110011011001011100111000000;
filter5[0][912] = 35'b11110100011111000001100111110000000;
filter5[0][913] = 35'b11111101110011000111100111100100000;
filter5[0][914] = 35'b00000001101100111011010100111100000;
filter5[0][915] = 35'b00000010010011110011111000000100000;
filter5[0][916] = 35'b11111111001010111111000001100011000;
filter5[0][917] = 35'b00000011101010000101100110011000000;
filter5[0][918] = 35'b00000000000110010011000001111111111;
filter5[0][919] = 35'b11111010011100001111110100111000000;
filter5[0][920] = 35'b11111011011010010000010011010000000;
filter5[0][921] = 35'b11111010100011111101001101010000000;
filter5[0][922] = 35'b00000010001100111111110100001100000;
filter5[0][923] = 35'b11111101100001111100100000000100000;
filter5[0][924] = 35'b00000000011001100011000101001001000;
filter5[0][925] = 35'b11111001101011100000011000110000000;
filter5[0][926] = 35'b00000011011011100011100111011100000;
filter5[0][927] = 35'b00000011100001110101000011001100000;
filter5[0][928] = 35'b00000001100100101111110001011000000;
filter5[0][929] = 35'b11111010011101110101101101111000000;
filter5[0][930] = 35'b00000001001011000011101001001010000;
filter5[0][931] = 35'b00000001101110100011011110010100000;
filter5[0][932] = 35'b00000011010010110111010110001000000;
filter5[0][933] = 35'b11111111111110010011000001100001111;
filter5[0][934] = 35'b11101101010110011111010100000000000;
filter5[0][935] = 35'b11110001011000011010110110100000000;
filter5[0][936] = 35'b11111101011001101011100000110100000;
filter5[0][937] = 35'b11111101011010000000011000001000000;
filter5[0][938] = 35'b11111101000010111101101001100000000;
filter5[0][939] = 35'b00000001100101101111010010010100000;
filter5[0][940] = 35'b11111111101111100001111001110101000;
filter5[0][941] = 35'b11111101000110101110100001010000000;
filter5[0][942] = 35'b11111101010100101101001100000000000;
filter5[0][943] = 35'b00000000110000111110100010001010000;
filter5[0][944] = 35'b11110110111010100101000011110000000;
filter5[0][945] = 35'b00000100010000010000111101101000000;
filter5[0][946] = 35'b00000000100011011010100011110001000;
filter5[0][947] = 35'b00000011000100111101110101111000000;
filter5[0][948] = 35'b11111101101100001101011011110100000;
filter5[0][949] = 35'b11111101011100000000111101110100000;
filter5[0][950] = 35'b00000001010110010100010111110100000;
filter5[0][951] = 35'b00000100110101011000101001000000000;
filter5[0][952] = 35'b11110111000111111111000010110000000;
filter5[0][953] = 35'b11111111111100100001100011010000111;
filter5[0][954] = 35'b00000010100110011110000011100100000;
filter5[0][955] = 35'b11111100100010000110011111111100000;
filter5[0][956] = 35'b11111011110001011101010101001000000;
filter5[0][957] = 35'b11101010011010010111011010100000000;
filter5[0][958] = 35'b11111011111000000100100110000000000;
filter5[0][959] = 35'b11111100100101111100011011011100000;
filter5[0][960] = 35'b00000000110000001010110101000011000;
filter5[0][961] = 35'b00000100111001001101001000110000000;
filter5[0][962] = 35'b00000000000011111101000101100101100;
filter5[0][963] = 35'b11111011100010001011110010011000000;
filter5[0][964] = 35'b00000011111010111101100010100000000;
filter5[0][965] = 35'b00000110110111100100101111001000000;
filter5[0][966] = 35'b00000110001110100011011101011000000;
filter5[0][967] = 35'b11111101000101001100000100100000000;
filter5[0][968] = 35'b00000010101110100101011111001100000;
filter5[0][969] = 35'b11111111011010101110100000000010000;
filter5[0][970] = 35'b11111110111001011000010101110110000;
filter5[0][971] = 35'b00000000111000111000010111010101000;
filter5[0][972] = 35'b11111111110011100101001110101111100;
filter5[0][973] = 35'b00000001010010001011010101001110000;
filter5[0][974] = 35'b11111110111101011011011011100010000;
filter5[0][975] = 35'b11111111000000010101001001110011000;
filter5[0][976] = 35'b11111100000000111111000100111100000;
filter5[0][977] = 35'b11111110101101110010100110100110000;
filter5[0][978] = 35'b11111111110101111001101001100101110;
filter5[0][979] = 35'b00000100000100101001101001100000000;
filter5[0][980] = 35'b11111111111001110011010010010010011;
filter5[0][981] = 35'b00000000010010000011101010110100000;
filter5[0][982] = 35'b00000001100111111110101100101000000;
filter5[0][983] = 35'b00000010111001001001001110000100000;
filter5[0][984] = 35'b11111010100010000100011110111000000;
filter5[0][985] = 35'b11110001111101111001100111010000000;
filter5[0][986] = 35'b00000010011001001010010110110100000;
filter5[0][987] = 35'b11111111011000110011110001101111000;
filter5[0][988] = 35'b00000010101100011110100011011100000;
filter5[0][989] = 35'b11111111100001000010000000101100000;
filter5[0][990] = 35'b00000000110101010101110010000111000;
filter5[0][991] = 35'b00000110001011100111011100000000000;
filter5[0][992] = 35'b11111010000100000101100010000000000;
filter5[0][993] = 35'b11111110011001001100110111100110000;
filter5[0][994] = 35'b11111100000011011101010110100000000;
filter5[0][995] = 35'b00000000101000010000000101100000000;
filter5[0][996] = 35'b00000100011010111001111000011000000;
filter5[0][997] = 35'b11111011111101011000000010100000000;
filter5[0][998] = 35'b11111111111111010110110110001011010;
filter5[0][999] = 35'b11111010000011111101110100111000000;
filter5[0][1000] = 35'b11110111110111100011100011000000000;
filter5[0][1001] = 35'b11111110111001001001111001000110000;
filter5[0][1002] = 35'b11111111110101000111000011010001010;
filter5[0][1003] = 35'b00000000011100010000011100101110000;
filter5[0][1004] = 35'b00000001100100111101011011010000000;
filter5[0][1005] = 35'b11111110011101111101001011000000000;
filter5[0][1006] = 35'b00000001001100100011110100011000000;
filter5[0][1007] = 35'b11111110100010111110001010100110000;
filter5[0][1008] = 35'b11111111001111110001001110101011000;
filter5[0][1009] = 35'b11111111010101000110001110101100000;
filter5[0][1010] = 35'b11111001010111101001100010000000000;
filter5[0][1011] = 35'b11111110000000000100101010010000000;
filter5[0][1012] = 35'b00000111100111011010001011010000000;
filter5[0][1013] = 35'b00000011010010110111000001101000000;
filter5[0][1014] = 35'b11111101010101001110111001111000000;
filter5[0][1015] = 35'b11111100101101111111101011111000000;
filter5[0][1016] = 35'b11111110110001001110111001011110000;
filter5[0][1017] = 35'b11111111110111010100110110111010110;
filter5[0][1018] = 35'b11111000001101001110100110100000000;
filter5[0][1019] = 35'b11110110111010011110100000100000000;
filter5[0][1020] = 35'b11101111110110010101001100000000000;
filter5[0][1021] = 35'b11111010001000001100000110011000000;
filter5[0][1022] = 35'b11110101111011100010101001110000000;
filter5[0][1023] = 35'b00000001111000110010110010110000000;
filter5[1][0] = 35'b00000000111101000110101100010011000;
filter5[1][1] = 35'b11111110010011101101001000111100000;
filter5[1][2] = 35'b00000000111111010000101110101010000;
filter5[1][3] = 35'b00000010000000100101000010000100000;
filter5[1][4] = 35'b00000101011101001001101110010000000;
filter5[1][5] = 35'b00000000000011110010110101100011001;
filter5[1][6] = 35'b11111111110011101001011111110000100;
filter5[1][7] = 35'b00000101011010110110011110101000000;
filter5[1][8] = 35'b11111100100001001110010101111000000;
filter5[1][9] = 35'b11111101111100110001001101100100000;
filter5[1][10] = 35'b00000000110111010100110011011111000;
filter5[1][11] = 35'b11110101101100100100111101000000000;
filter5[1][12] = 35'b00000110111101110100010010100000000;
filter5[1][13] = 35'b11111101010011100111000110100000000;
filter5[1][14] = 35'b11111110000010001110101110011110000;
filter5[1][15] = 35'b00000100101110010011010011100000000;
filter5[1][16] = 35'b00000000100110001000010010100010000;
filter5[1][17] = 35'b00000000100111001000011100000100000;
filter5[1][18] = 35'b11111110110000011111111000111110000;
filter5[1][19] = 35'b11111101010000000101001001011100000;
filter5[1][20] = 35'b11111101100101110011010100000000000;
filter5[1][21] = 35'b11111111101100001101000100010111100;
filter5[1][22] = 35'b00000001101010111111010001011110000;
filter5[1][23] = 35'b00000111110100110101100001010000000;
filter5[1][24] = 35'b00000010111011111110111100010000000;
filter5[1][25] = 35'b00000010000100010000110000101100000;
filter5[1][26] = 35'b11111111010101001111101110000011000;
filter5[1][27] = 35'b11111010110000101111100101110000000;
filter5[1][28] = 35'b00000000011000001110100101100010100;
filter5[1][29] = 35'b11111111000011011010111001000010000;
filter5[1][30] = 35'b00000011100110110110010100000100000;
filter5[1][31] = 35'b11111011101001111100010011000000000;
filter5[1][32] = 35'b00000001011111110011100100101000000;
filter5[1][33] = 35'b00000100001111000101010010101000000;
filter5[1][34] = 35'b00000011101001100101110011011000000;
filter5[1][35] = 35'b00000000110110100111110011010011000;
filter5[1][36] = 35'b00000011110000110000001001000000000;
filter5[1][37] = 35'b11111001100111100011010111000000000;
filter5[1][38] = 35'b00000010111011011110100000010100000;
filter5[1][39] = 35'b11111010111000000111000110000000000;
filter5[1][40] = 35'b11111110110000111100001101001110000;
filter5[1][41] = 35'b11111100100011010011010010101000000;
filter5[1][42] = 35'b00000001000010101100110010100100000;
filter5[1][43] = 35'b00000000000010110100010001101100001;
filter5[1][44] = 35'b11111101111011111010111001001100000;
filter5[1][45] = 35'b00000010101010000000000111101100000;
filter5[1][46] = 35'b11111111110110111111101110100001100;
filter5[1][47] = 35'b11111010101001000001101010010000000;
filter5[1][48] = 35'b11110111011101001001101101000000000;
filter5[1][49] = 35'b00000001001011111011101101001100000;
filter5[1][50] = 35'b00000001010011001011101101000010000;
filter5[1][51] = 35'b11111101110000010110001101111100000;
filter5[1][52] = 35'b00000001101111101001111001011000000;
filter5[1][53] = 35'b11111111000101010010111110100000000;
filter5[1][54] = 35'b00000000011101000000001101100110000;
filter5[1][55] = 35'b11111100111111000001010110001100000;
filter5[1][56] = 35'b00000000000101110011000110110001110;
filter5[1][57] = 35'b00000011000011000011000110110100000;
filter5[1][58] = 35'b00000001011000100011011100001000000;
filter5[1][59] = 35'b11111100000010111011110100101000000;
filter5[1][60] = 35'b00000001000001111000110101010110000;
filter5[1][61] = 35'b11111111101011100100100011010110000;
filter5[1][62] = 35'b00000011010110100110001011110000000;
filter5[1][63] = 35'b11111100100011111101011000010100000;
filter5[1][64] = 35'b11111101110100110100000100100100000;
filter5[1][65] = 35'b00000001000111101100001111100110000;
filter5[1][66] = 35'b00000001100100100101100110111010000;
filter5[1][67] = 35'b11111110100101110110101110101110000;
filter5[1][68] = 35'b00000000010011110111001010110010100;
filter5[1][69] = 35'b11111111111110011100100110001011100;
filter5[1][70] = 35'b00000001110001001101111100101100000;
filter5[1][71] = 35'b00000001011001110111010101011110000;
filter5[1][72] = 35'b11111101111011100110010100101100000;
filter5[1][73] = 35'b11111111101010001111101010011111000;
filter5[1][74] = 35'b00000010011000111010100011001100000;
filter5[1][75] = 35'b11111111101100111001000010010000000;
filter5[1][76] = 35'b11111111000101100000100100000100000;
filter5[1][77] = 35'b11111110101110101011111011110100000;
filter5[1][78] = 35'b11111101001100100000100011001000000;
filter5[1][79] = 35'b11111101110110100100110010100000000;
filter5[1][80] = 35'b00000000111000000000011001101110000;
filter5[1][81] = 35'b00000001100000000101011101111110000;
filter5[1][82] = 35'b00000000111111011101101101001111000;
filter5[1][83] = 35'b11111110000000000101000001101110000;
filter5[1][84] = 35'b11111110101011100011111000011100000;
filter5[1][85] = 35'b11111110011000000100001101101110000;
filter5[1][86] = 35'b11111110111010000011110100010100000;
filter5[1][87] = 35'b00000010011100101100001011111000000;
filter5[1][88] = 35'b00000100010111000001100101011000000;
filter5[1][89] = 35'b00000010101000100000110100001100000;
filter5[1][90] = 35'b00000001100100010010100011011000000;
filter5[1][91] = 35'b11111101100001100110011011111000000;
filter5[1][92] = 35'b00000000110111111000001101010111000;
filter5[1][93] = 35'b11111111000011010110110001010100000;
filter5[1][94] = 35'b00000100101110110110001000000000000;
filter5[1][95] = 35'b11111101001110101111111010001000000;
filter5[1][96] = 35'b11111101100011011010110000111100000;
filter5[1][97] = 35'b00000100111000101000011011110000000;
filter5[1][98] = 35'b00000011110111110111111100101100000;
filter5[1][99] = 35'b00000000011000011100010100000010000;
filter5[1][100] = 35'b00000011111101010011010001010100000;
filter5[1][101] = 35'b11111100101010001111110100000100000;
filter5[1][102] = 35'b11111100011101101100000011111000000;
filter5[1][103] = 35'b00000001010111001101110000110010000;
filter5[1][104] = 35'b00000000001000011011010100100001010;
filter5[1][105] = 35'b00000001011000110100000011001110000;
filter5[1][106] = 35'b00000000101011000100001011100000000;
filter5[1][107] = 35'b11111011011001011000111100000000000;
filter5[1][108] = 35'b00000000000111001001011001011000100;
filter5[1][109] = 35'b00000001100001100111110111111010000;
filter5[1][110] = 35'b00000000101011001100010101000110000;
filter5[1][111] = 35'b11111110100100111011101000010010000;
filter5[1][112] = 35'b11111101100011101110110101011100000;
filter5[1][113] = 35'b11111111001111100011110011101000000;
filter5[1][114] = 35'b11111101110001010010101100000000000;
filter5[1][115] = 35'b11111110000101001010101010000000000;
filter5[1][116] = 35'b00000011011011100010101010010100000;
filter5[1][117] = 35'b11111110110010110111100100101100000;
filter5[1][118] = 35'b00000000001110010111100011000010000;
filter5[1][119] = 35'b00000000111011011110100101101101000;
filter5[1][120] = 35'b00000010011111111010011100010000000;
filter5[1][121] = 35'b00000001110010001110100001011100000;
filter5[1][122] = 35'b11111101010001100001101110100000000;
filter5[1][123] = 35'b11111100110011010110111101001000000;
filter5[1][124] = 35'b00000000100011001010000111100110000;
filter5[1][125] = 35'b00000000110101001101010101010110000;
filter5[1][126] = 35'b11111101000110001110110010100000000;
filter5[1][127] = 35'b11111100110110000010011101000000000;
filter5[1][128] = 35'b11110100110010001100111101110000000;
filter5[1][129] = 35'b11111100000011111100011100111100000;
filter5[1][130] = 35'b11111011000101100101001000011000000;
filter5[1][131] = 35'b11110001111011110011000010100000000;
filter5[1][132] = 35'b00000000011010011010101001110001100;
filter5[1][133] = 35'b00000010111110011101001110110000000;
filter5[1][134] = 35'b00000010110111000000110110110100000;
filter5[1][135] = 35'b00000011100000000101001010001000000;
filter5[1][136] = 35'b11111011100111100100110010111000000;
filter5[1][137] = 35'b11111101100101001110100010110100000;
filter5[1][138] = 35'b00000101101000100101011010000000000;
filter5[1][139] = 35'b00000000100100101111111100111011000;
filter5[1][140] = 35'b11111110011101011010000010001000000;
filter5[1][141] = 35'b11101010111000010000011001000000000;
filter5[1][142] = 35'b11110011111101010110010011000000000;
filter5[1][143] = 35'b11111100111001010100100100101100000;
filter5[1][144] = 35'b00000100001101011101010111111000000;
filter5[1][145] = 35'b00000001000111011011110100001100000;
filter5[1][146] = 35'b00000000110010111111000001001000000;
filter5[1][147] = 35'b11111111110111001001100010110011000;
filter5[1][148] = 35'b11111111101001011010110111100101000;
filter5[1][149] = 35'b00000010100010000100001011101000000;
filter5[1][150] = 35'b11110001110011010011011111110000000;
filter5[1][151] = 35'b00000000010110100111110011110110100;
filter5[1][152] = 35'b00000111000110111001100110111000000;
filter5[1][153] = 35'b00000010101111010010100111000100000;
filter5[1][154] = 35'b00000101000110100111010011001000000;
filter5[1][155] = 35'b00000010000101011011000110100000000;
filter5[1][156] = 35'b11111100000100100010100001110000000;
filter5[1][157] = 35'b11111001110001110110011111011000000;
filter5[1][158] = 35'b11111110110100010111001101011010000;
filter5[1][159] = 35'b11110110000100100111011011110000000;
filter5[1][160] = 35'b00001001000010101001111000100000000;
filter5[1][161] = 35'b00001110101001101110110110010000000;
filter5[1][162] = 35'b00000100000011000011101101010000000;
filter5[1][163] = 35'b00000010101000000000010101001000000;
filter5[1][164] = 35'b11111111100100111000010001011010100;
filter5[1][165] = 35'b11110110110011010110011000010000000;
filter5[1][166] = 35'b11111100011111100001101011000100000;
filter5[1][167] = 35'b11111001110101110101111000001000000;
filter5[1][168] = 35'b00000001000011110110011101000010000;
filter5[1][169] = 35'b11111111011100100010101011001111000;
filter5[1][170] = 35'b11111111110000000011010100011011010;
filter5[1][171] = 35'b00000001011010110000001110000110000;
filter5[1][172] = 35'b11111011111111101111001001101000000;
filter5[1][173] = 35'b11111111001110000011001101001001000;
filter5[1][174] = 35'b11110010010000111000000110100000000;
filter5[1][175] = 35'b11110010001010001110110101100000000;
filter5[1][176] = 35'b11111100101110110100111100100100000;
filter5[1][177] = 35'b11101101111010111100110001100000000;
filter5[1][178] = 35'b11110010101111011000011101110000000;
filter5[1][179] = 35'b11111011010001001000111011011000000;
filter5[1][180] = 35'b11111110010000101010100000011100000;
filter5[1][181] = 35'b00000000101001010101000000001100000;
filter5[1][182] = 35'b11111101110101010111100110111000000;
filter5[1][183] = 35'b11110101100011111011101111000000000;
filter5[1][184] = 35'b11110010001110001011100011010000000;
filter5[1][185] = 35'b11111011010010001011110010100000000;
filter5[1][186] = 35'b11111100010110111111101101001000000;
filter5[1][187] = 35'b11110011110000011011011110100000000;
filter5[1][188] = 35'b11111011010001011000100111101000000;
filter5[1][189] = 35'b11111111111001100111011100110001001;
filter5[1][190] = 35'b11110000010100010001001000000000000;
filter5[1][191] = 35'b11110010111000000000001101110000000;
filter5[1][192] = 35'b11110111001111011000101101100000000;
filter5[1][193] = 35'b11101110011000101111001111000000000;
filter5[1][194] = 35'b11111100111000000011000100000100000;
filter5[1][195] = 35'b00000001001000111100101110100010000;
filter5[1][196] = 35'b11111010010101011111101000010000000;
filter5[1][197] = 35'b11111110011011110010001101110000000;
filter5[1][198] = 35'b11111111100100110001000010110010100;
filter5[1][199] = 35'b00001000101110100010000101110000000;
filter5[1][200] = 35'b11111010100100111101000100111000000;
filter5[1][201] = 35'b11110110110010101010110001010000000;
filter5[1][202] = 35'b11111110100110011101100101000110000;
filter5[1][203] = 35'b11111001111000010010000110100000000;
filter5[1][204] = 35'b11110101100001001000011010010000000;
filter5[1][205] = 35'b11110110010011010010011010000000000;
filter5[1][206] = 35'b11111100101000001011101011100000000;
filter5[1][207] = 35'b11111011111100111110101011010000000;
filter5[1][208] = 35'b11110101100110111001101110010000000;
filter5[1][209] = 35'b00000011000001010111101100011100000;
filter5[1][210] = 35'b11111110101101010111011110001000000;
filter5[1][211] = 35'b11111110001011100010011000101000000;
filter5[1][212] = 35'b00000010000100111010111111101000000;
filter5[1][213] = 35'b11111111010000011100011110101000000;
filter5[1][214] = 35'b11111010010001000011001011111000000;
filter5[1][215] = 35'b00000000000011010101001111100100101;
filter5[1][216] = 35'b11110111001000110101010100110000000;
filter5[1][217] = 35'b00000101010001111110011000011000000;
filter5[1][218] = 35'b11111110101001010111000000100110000;
filter5[1][219] = 35'b11111110011010001101001001001000000;
filter5[1][220] = 35'b00000000001010010011000000001100100;
filter5[1][221] = 35'b11111110101110000000000101001000000;
filter5[1][222] = 35'b11110001010011111000101110000000000;
filter5[1][223] = 35'b11111110110110100111011100000110000;
filter5[1][224] = 35'b11111011101100110000000111100000000;
filter5[1][225] = 35'b11111001101111100011100100011000000;
filter5[1][226] = 35'b00000110001111010101110111010000000;
filter5[1][227] = 35'b11111110111110110000011010011000000;
filter5[1][228] = 35'b00000011001101001000101010111000000;
filter5[1][229] = 35'b00000010100001100011011100011000000;
filter5[1][230] = 35'b11111100001000111110000000000000000;
filter5[1][231] = 35'b00000100000111110001110100010000000;
filter5[1][232] = 35'b11111000110000001110101100010000000;
filter5[1][233] = 35'b11111111011100110000101001101000000;
filter5[1][234] = 35'b00000011110001010001110110000000000;
filter5[1][235] = 35'b00000001111010011001011001010100000;
filter5[1][236] = 35'b11111010101011101010101011110000000;
filter5[1][237] = 35'b00000001001101111111000110000010000;
filter5[1][238] = 35'b00000000011101110110010110001111000;
filter5[1][239] = 35'b11111110100101001111100101001010000;
filter5[1][240] = 35'b11110111010010100001110101100000000;
filter5[1][241] = 35'b11111110000101100010011001011110000;
filter5[1][242] = 35'b00000001000111010011100011000100000;
filter5[1][243] = 35'b11111011101011111110101010100000000;
filter5[1][244] = 35'b11111110001100110010011000000110000;
filter5[1][245] = 35'b11111110010001110010011111110000000;
filter5[1][246] = 35'b11111111010100010000111000111100000;
filter5[1][247] = 35'b11111110110010001111001000011110000;
filter5[1][248] = 35'b11110101000101010111110110110000000;
filter5[1][249] = 35'b11111110000011011100100100100100000;
filter5[1][250] = 35'b11111101001011010111011111101100000;
filter5[1][251] = 35'b11111110001011001101000110011010000;
filter5[1][252] = 35'b11111100110010011010010010001100000;
filter5[1][253] = 35'b00000010101000100011000001001000000;
filter5[1][254] = 35'b00000010111010110011001000011100000;
filter5[1][255] = 35'b11111000010100110000000101110000000;
filter5[1][256] = 35'b11111000011101101001010000111000000;
filter5[1][257] = 35'b00000000011010100010100011011111000;
filter5[1][258] = 35'b11111011001110000001010101011000000;
filter5[1][259] = 35'b11111001010110111110111000010000000;
filter5[1][260] = 35'b11111101011101111011111100101000000;
filter5[1][261] = 35'b11111100101110100000100010001100000;
filter5[1][262] = 35'b11111111011110001101000101000011000;
filter5[1][263] = 35'b00000000011000001000000100010100100;
filter5[1][264] = 35'b11111010001001111101011001111000000;
filter5[1][265] = 35'b11110100010000010111100010100000000;
filter5[1][266] = 35'b11111011100101010111111111011000000;
filter5[1][267] = 35'b11110111110001101101001000110000000;
filter5[1][268] = 35'b11110110000101000010110000000000000;
filter5[1][269] = 35'b11111111011111000111001101011011000;
filter5[1][270] = 35'b11111101111101011101101111000100000;
filter5[1][271] = 35'b11111111001010101110100010101100000;
filter5[1][272] = 35'b00000001001001110010011100110010000;
filter5[1][273] = 35'b00000011000001101100001000000000000;
filter5[1][274] = 35'b11111101100001100001101100110000000;
filter5[1][275] = 35'b11111100111000011100101101011000000;
filter5[1][276] = 35'b00000001000010000111101100101100000;
filter5[1][277] = 35'b11111011100011101011100010110000000;
filter5[1][278] = 35'b11111100101001011110000111001000000;
filter5[1][279] = 35'b11111110110100111010100100010100000;
filter5[1][280] = 35'b11111100100100001001001111101100000;
filter5[1][281] = 35'b00000001000110110101010111011010000;
filter5[1][282] = 35'b00000010100011011110010111101000000;
filter5[1][283] = 35'b00000000000101110101100111000101100;
filter5[1][284] = 35'b00000000101000100001001011001111000;
filter5[1][285] = 35'b11111100101001100011011000110100000;
filter5[1][286] = 35'b11111101000001110011111001010000000;
filter5[1][287] = 35'b11111101000100111010011110011000000;
filter5[1][288] = 35'b11111101000111011111000001101000000;
filter5[1][289] = 35'b11111110101001011001001101111100000;
filter5[1][290] = 35'b00000010111110000000100011000000000;
filter5[1][291] = 35'b11111111100001110101100101001010000;
filter5[1][292] = 35'b11111110001101111001110110001010000;
filter5[1][293] = 35'b11111010110111000010000001100000000;
filter5[1][294] = 35'b11111100100111101110011100101100000;
filter5[1][295] = 35'b11111011101101100011111101001000000;
filter5[1][296] = 35'b00000100011011011110000101000000000;
filter5[1][297] = 35'b11111000010001011111111000000000000;
filter5[1][298] = 35'b00000001101001110110100100101100000;
filter5[1][299] = 35'b11111100011100100000100110010000000;
filter5[1][300] = 35'b11111110001000000001011000111010000;
filter5[1][301] = 35'b11111101011001111011000001100000000;
filter5[1][302] = 35'b11111010011011101000000100101000000;
filter5[1][303] = 35'b11111011110110111001100111111000000;
filter5[1][304] = 35'b11110100000010010010111111000000000;
filter5[1][305] = 35'b00000001000110011100110011000110000;
filter5[1][306] = 35'b00000010110010001001011010101100000;
filter5[1][307] = 35'b11111100111010101101010110100100000;
filter5[1][308] = 35'b11111011011010100001100101101000000;
filter5[1][309] = 35'b11111111111001110001000110111000010;
filter5[1][310] = 35'b11111001101111010011011011100000000;
filter5[1][311] = 35'b11111101000000010001111110111100000;
filter5[1][312] = 35'b11110001100100010101100110100000000;
filter5[1][313] = 35'b11110110101100000111100010000000000;
filter5[1][314] = 35'b11111001010111010100111110111000000;
filter5[1][315] = 35'b00000000101011011101001000101011000;
filter5[1][316] = 35'b11111111110011010101000010001111110;
filter5[1][317] = 35'b00000101000010001010110110011000000;
filter5[1][318] = 35'b11111000100101011101110111100000000;
filter5[1][319] = 35'b11111010011111111011001011111000000;
filter5[1][320] = 35'b00000010001011110001001001110000000;
filter5[1][321] = 35'b11111111101100100010110010110001100;
filter5[1][322] = 35'b11111111000100011100111001010100000;
filter5[1][323] = 35'b11111111111110111110100111100000001;
filter5[1][324] = 35'b11111111100001011011001111010011100;
filter5[1][325] = 35'b00000010010111101001101001100100000;
filter5[1][326] = 35'b00000010111010000101011100110000000;
filter5[1][327] = 35'b00001000011010001010111111010000000;
filter5[1][328] = 35'b11111010100001001100111000010000000;
filter5[1][329] = 35'b11111110010111010010011010100100000;
filter5[1][330] = 35'b00000010110000001101001011010100000;
filter5[1][331] = 35'b00000000011011010111110101111010100;
filter5[1][332] = 35'b11111111011001111000101101001101000;
filter5[1][333] = 35'b11110001111101001000001100100000000;
filter5[1][334] = 35'b00000001101010010100101000011110000;
filter5[1][335] = 35'b00000011101010100010011011111100000;
filter5[1][336] = 35'b00000001110000010000001100001110000;
filter5[1][337] = 35'b00000001011001000000000001101110000;
filter5[1][338] = 35'b11111110000110010100011110001100000;
filter5[1][339] = 35'b11111100101110111110000010010100000;
filter5[1][340] = 35'b11111101110011000101100100001000000;
filter5[1][341] = 35'b11111110111100110111010001011000000;
filter5[1][342] = 35'b11111100111000100100000101110000000;
filter5[1][343] = 35'b00000001110001001000010011101110000;
filter5[1][344] = 35'b11111111011111101111011100000001000;
filter5[1][345] = 35'b00000001100111111010010100001000000;
filter5[1][346] = 35'b00000000000000111011101100010111100;
filter5[1][347] = 35'b00000010000100011110100100101100000;
filter5[1][348] = 35'b00000101010111001101111001011000000;
filter5[1][349] = 35'b00000001011110000110110011000000000;
filter5[1][350] = 35'b11111110101001001111110000100100000;
filter5[1][351] = 35'b11111101100101101101100001111000000;
filter5[1][352] = 35'b00000000010110100110010110101100100;
filter5[1][353] = 35'b11111011101011011011111110001000000;
filter5[1][354] = 35'b00000100100001011010001110010000000;
filter5[1][355] = 35'b00000000000001101000110000101011101;
filter5[1][356] = 35'b00000000010000110110101000000100100;
filter5[1][357] = 35'b11111100000000011011111110011100000;
filter5[1][358] = 35'b00000010001100100101111000011100000;
filter5[1][359] = 35'b11111001111101010000010110111000000;
filter5[1][360] = 35'b11111111011110101000000001100011000;
filter5[1][361] = 35'b11111111101101110101111011001101100;
filter5[1][362] = 35'b11111111011000001010010111011011000;
filter5[1][363] = 35'b11111110110110001110010000111010000;
filter5[1][364] = 35'b11111111010001101001101001111011000;
filter5[1][365] = 35'b11111110101001100011000100100010000;
filter5[1][366] = 35'b11111101110001101110110100001000000;
filter5[1][367] = 35'b11111110111010111110110110101110000;
filter5[1][368] = 35'b11111101001010001101110110101100000;
filter5[1][369] = 35'b11111101100000111100000000010000000;
filter5[1][370] = 35'b11111110011001100010010110101010000;
filter5[1][371] = 35'b11111111110111001011101101000110110;
filter5[1][372] = 35'b11111011001110110101001101000000000;
filter5[1][373] = 35'b11111111011011010001000100010110000;
filter5[1][374] = 35'b00000001101000000100111101111010000;
filter5[1][375] = 35'b11111111010010110000101010010001000;
filter5[1][376] = 35'b11111000100010010010110011011000000;
filter5[1][377] = 35'b11111111101001111001100000111011100;
filter5[1][378] = 35'b11111111111111000001111001111000110;
filter5[1][379] = 35'b11111101010100001111001111001000000;
filter5[1][380] = 35'b00000010110011101100001010011000000;
filter5[1][381] = 35'b00000011010110001010000101111100000;
filter5[1][382] = 35'b00000010001001000001101010000100000;
filter5[1][383] = 35'b11111100000001011000001101101000000;
filter5[1][384] = 35'b00000010111110101101111111011000000;
filter5[1][385] = 35'b00000000110110001010010010111001000;
filter5[1][386] = 35'b11111111000110011101110110001100000;
filter5[1][387] = 35'b00000000111101011101000111111111000;
filter5[1][388] = 35'b11111101010101001100001010100000000;
filter5[1][389] = 35'b11111110101010001101000011010000000;
filter5[1][390] = 35'b11111101010101110001010011000000000;
filter5[1][391] = 35'b11111101011000011000000100001100000;
filter5[1][392] = 35'b11111100111001101110001110000100000;
filter5[1][393] = 35'b11111111010101011110000010000000000;
filter5[1][394] = 35'b11111110000000111101111001100010000;
filter5[1][395] = 35'b11111111101100001000100011000100100;
filter5[1][396] = 35'b00000001110110101110001000000100000;
filter5[1][397] = 35'b00000001110011001110010010001100000;
filter5[1][398] = 35'b00000000010111000100010111010111000;
filter5[1][399] = 35'b11111111110001010101100011000001110;
filter5[1][400] = 35'b00000011101101010101110101101000000;
filter5[1][401] = 35'b00000010100000010000101000001100000;
filter5[1][402] = 35'b11111110100000101000000011100000000;
filter5[1][403] = 35'b11111100010011010000001001000100000;
filter5[1][404] = 35'b11111111001100111110010111111001000;
filter5[1][405] = 35'b00000000100011100011101110100100000;
filter5[1][406] = 35'b11111111111111010010000101111010010;
filter5[1][407] = 35'b11111111010001001110001111010111000;
filter5[1][408] = 35'b00000000110010100011110010000001000;
filter5[1][409] = 35'b00000010001100001110101010101000000;
filter5[1][410] = 35'b00000000011101110111001111011001000;
filter5[1][411] = 35'b00000010011000111111010101101000000;
filter5[1][412] = 35'b00000001111000000011011000100110000;
filter5[1][413] = 35'b11111111110111010111011101011000010;
filter5[1][414] = 35'b00000100011101111111110001110000000;
filter5[1][415] = 35'b00000011101001001101000011000000000;
filter5[1][416] = 35'b11111110011111010100011111110000000;
filter5[1][417] = 35'b11111101001111101111000110101000000;
filter5[1][418] = 35'b11111101110110100100101100100100000;
filter5[1][419] = 35'b00000000111111110001010011110110000;
filter5[1][420] = 35'b11111110011100100010010110001100000;
filter5[1][421] = 35'b00000101100111000111000001110000000;
filter5[1][422] = 35'b11111011011010101001100111001000000;
filter5[1][423] = 35'b00000001000111001111000111110000000;
filter5[1][424] = 35'b00000001000100101001001101101110000;
filter5[1][425] = 35'b00000011100001000110000111011000000;
filter5[1][426] = 35'b11111110110101110011111010111000000;
filter5[1][427] = 35'b00000011101110111011001100110100000;
filter5[1][428] = 35'b00000000100011111111011100111110000;
filter5[1][429] = 35'b11111101100011000010100101111000000;
filter5[1][430] = 35'b11111101000000000110000110011000000;
filter5[1][431] = 35'b11111110100001001001001010010110000;
filter5[1][432] = 35'b00000000101111011101001001111001000;
filter5[1][433] = 35'b00000001101011110011100001110110000;
filter5[1][434] = 35'b11111111110010101000010111010101110;
filter5[1][435] = 35'b11111111011011011101011111110001000;
filter5[1][436] = 35'b00000000011010100000101011111101100;
filter5[1][437] = 35'b00000000000101011000000010000000000;
filter5[1][438] = 35'b11111110111010101100011000010000000;
filter5[1][439] = 35'b00000000111000010011110100101111000;
filter5[1][440] = 35'b11111101111011000101111010100100000;
filter5[1][441] = 35'b11111110100000000111101000110010000;
filter5[1][442] = 35'b00000000010010110000101001111000000;
filter5[1][443] = 35'b11111110111010010011001000110010000;
filter5[1][444] = 35'b11111101001001001011100101100000000;
filter5[1][445] = 35'b00000000010001000011111001000100000;
filter5[1][446] = 35'b00000010100000100001011010101000000;
filter5[1][447] = 35'b00000100111101100110010010100000000;
filter5[1][448] = 35'b00000101000011010101000010100000000;
filter5[1][449] = 35'b00000000111100001001110011010101000;
filter5[1][450] = 35'b00000100010100101010000111000000000;
filter5[1][451] = 35'b00000101111000011110111110001000000;
filter5[1][452] = 35'b11111011110111000001011011010000000;
filter5[1][453] = 35'b11111111001010001001100011010010000;
filter5[1][454] = 35'b11111010111101000010000111100000000;
filter5[1][455] = 35'b11111010000001100110111110000000000;
filter5[1][456] = 35'b00000001101011101101011111001100000;
filter5[1][457] = 35'b11111100110000010101100010010100000;
filter5[1][458] = 35'b11111100111001101101011011100100000;
filter5[1][459] = 35'b11111111100111110100010111101110000;
filter5[1][460] = 35'b00000011000111110111110111101100000;
filter5[1][461] = 35'b00000100101100100101000000110000000;
filter5[1][462] = 35'b11111011100100010001100101110000000;
filter5[1][463] = 35'b00000011110000101011101101110100000;
filter5[1][464] = 35'b00000110001001010111011010001000000;
filter5[1][465] = 35'b11111101111101010001010001111000000;
filter5[1][466] = 35'b11101010110111110000111111100000000;
filter5[1][467] = 35'b11111110010101011001100000110010000;
filter5[1][468] = 35'b11111110100101011101100110101110000;
filter5[1][469] = 35'b11111011100010011110000000001000000;
filter5[1][470] = 35'b11111101100101001010010001001100000;
filter5[1][471] = 35'b00000001001011100010011100100010000;
filter5[1][472] = 35'b00010000110111000010110110100000000;
filter5[1][473] = 35'b00000110001100100110111001100000000;
filter5[1][474] = 35'b00000010010010011111000010011100000;
filter5[1][475] = 35'b00000101110101100101111010110000000;
filter5[1][476] = 35'b11111111011100011110111010000001000;
filter5[1][477] = 35'b11111100100010010101011001001000000;
filter5[1][478] = 35'b11111000010110111101011011110000000;
filter5[1][479] = 35'b00000011001011011111000011111100000;
filter5[1][480] = 35'b00001001000001011101100101110000000;
filter5[1][481] = 35'b00010111001101000010001111000000000;
filter5[1][482] = 35'b00001000110001110110101000010000000;
filter5[1][483] = 35'b00000010011101110001110001011100000;
filter5[1][484] = 35'b00000000111111000001000011100011000;
filter5[1][485] = 35'b00000010010001100101110011001000000;
filter5[1][486] = 35'b11111010111010010001110000000000000;
filter5[1][487] = 35'b00000001100100010000111111110000000;
filter5[1][488] = 35'b11111101111111011001001010001100000;
filter5[1][489] = 35'b00000101101001010010001000101000000;
filter5[1][490] = 35'b00000010000010010101010001110000000;
filter5[1][491] = 35'b00000011110110011100111010110000000;
filter5[1][492] = 35'b00000000101110101101010001001000000;
filter5[1][493] = 35'b11111101011100110010100000000100000;
filter5[1][494] = 35'b11111100101111110111000101110100000;
filter5[1][495] = 35'b11111011001100001010100000110000000;
filter5[1][496] = 35'b11111111110101000111010001000111000;
filter5[1][497] = 35'b00000000100111100101000010101100000;
filter5[1][498] = 35'b11111111101000001101001010100111100;
filter5[1][499] = 35'b11111101111011110110111011000100000;
filter5[1][500] = 35'b11110111110101110110100100100000000;
filter5[1][501] = 35'b11111100111011010111110101011100000;
filter5[1][502] = 35'b00000000011010010100100001100010100;
filter5[1][503] = 35'b11111101101110000111110100111000000;
filter5[1][504] = 35'b11111000111101111111001111011000000;
filter5[1][505] = 35'b00000100110000011111001110000000000;
filter5[1][506] = 35'b00000000011011000110000010100101000;
filter5[1][507] = 35'b00000000010100001011010011101100000;
filter5[1][508] = 35'b11111100011010110000010011111000000;
filter5[1][509] = 35'b11110111101111100101000011100000000;
filter5[1][510] = 35'b11111110001000010001010101000010000;
filter5[1][511] = 35'b00000000101000001001011100000110000;
filter5[1][512] = 35'b00000000110001101100110111100001000;
filter5[1][513] = 35'b00000000001010101011110010000010010;
filter5[1][514] = 35'b00000000000100101001111001101001011;
filter5[1][515] = 35'b11111111110110100010100101001011010;
filter5[1][516] = 35'b11111110011110001101101000011000000;
filter5[1][517] = 35'b00000010001010111011000010110000000;
filter5[1][518] = 35'b11111110111100111000010101011000000;
filter5[1][519] = 35'b00000011111010111001100111010100000;
filter5[1][520] = 35'b00000000010001110010101110000100000;
filter5[1][521] = 35'b00000001010000010011000011001110000;
filter5[1][522] = 35'b11111110111011010010010010111100000;
filter5[1][523] = 35'b11111101001011111110001001011000000;
filter5[1][524] = 35'b00000011110010100101101110010100000;
filter5[1][525] = 35'b11111101000010101100011001100100000;
filter5[1][526] = 35'b11111111111011101000111101110110000;
filter5[1][527] = 35'b00000010110010110111001011010000000;
filter5[1][528] = 35'b00000011011010001110010001110000000;
filter5[1][529] = 35'b00000011100100011000101111011100000;
filter5[1][530] = 35'b11111111110001010010111001011011010;
filter5[1][531] = 35'b11111100111011011000101100111000000;
filter5[1][532] = 35'b11111110100101001010000010000110000;
filter5[1][533] = 35'b11111101000100111001100100001000000;
filter5[1][534] = 35'b00000010000101110110100011010100000;
filter5[1][535] = 35'b00000001011101101001001011001100000;
filter5[1][536] = 35'b00000010100011110000101101000100000;
filter5[1][537] = 35'b11111110111000110010010101111100000;
filter5[1][538] = 35'b11111111110111000111110110110010000;
filter5[1][539] = 35'b11111111010010101101010111101001000;
filter5[1][540] = 35'b00000010010001010011000111011100000;
filter5[1][541] = 35'b00000000000110110011010111011011001;
filter5[1][542] = 35'b11111110111010110011000110111110000;
filter5[1][543] = 35'b00000100010011101011111011001000000;
filter5[1][544] = 35'b00000011011111100010000001010100000;
filter5[1][545] = 35'b00000100101100000110011100111000000;
filter5[1][546] = 35'b00000000101100001100111011000111000;
filter5[1][547] = 35'b00000000001001011010101000110110110;
filter5[1][548] = 35'b00000010101001000111010111101000000;
filter5[1][549] = 35'b11111100110101111001110000101100000;
filter5[1][550] = 35'b00000000011000110010100010010100100;
filter5[1][551] = 35'b11111100111101010111101100011100000;
filter5[1][552] = 35'b00000000001010100100101111001101110;
filter5[1][553] = 35'b11111111010011001001001000001111000;
filter5[1][554] = 35'b00000100110001101001000110111000000;
filter5[1][555] = 35'b11111110110000010001100000110100000;
filter5[1][556] = 35'b11111111110010100001011010000001100;
filter5[1][557] = 35'b11111101010111010011100100110000000;
filter5[1][558] = 35'b11111101111101010101011000000000000;
filter5[1][559] = 35'b11111110001001011111111101111000000;
filter5[1][560] = 35'b11111101100101111001101000011100000;
filter5[1][561] = 35'b11111111100100110001101010100011100;
filter5[1][562] = 35'b11111011101111101100101001011000000;
filter5[1][563] = 35'b11111100101011011010000101000000000;
filter5[1][564] = 35'b11111110011000110010110000111110000;
filter5[1][565] = 35'b11111110111111001010101100010100000;
filter5[1][566] = 35'b00000010011000011101110001111000000;
filter5[1][567] = 35'b00000010101101010111001110010000000;
filter5[1][568] = 35'b11111011111100011011110011111000000;
filter5[1][569] = 35'b00000010010111010111111010001000000;
filter5[1][570] = 35'b00000100000000111000110011100000000;
filter5[1][571] = 35'b00000000110000010101101010000010000;
filter5[1][572] = 35'b11111110000111011010110111111100000;
filter5[1][573] = 35'b00000011100000011000001110000000000;
filter5[1][574] = 35'b00000001100101001010000110011010000;
filter5[1][575] = 35'b00000001101010001001010010000100000;
filter5[1][576] = 35'b11111101110000011011010101001000000;
filter5[1][577] = 35'b11111111101100100101101010000111000;
filter5[1][578] = 35'b00000000001110011110100110010111110;
filter5[1][579] = 35'b00000010010001111010100111100000000;
filter5[1][580] = 35'b11111011100010011000000001010000000;
filter5[1][581] = 35'b11111101001110110111100101111100000;
filter5[1][582] = 35'b11111100010100001100000001101000000;
filter5[1][583] = 35'b00000010111101001000011001100000000;
filter5[1][584] = 35'b00000000100001111101001011000011000;
filter5[1][585] = 35'b00000000111001011111010110100100000;
filter5[1][586] = 35'b11111010000011011000011100010000000;
filter5[1][587] = 35'b11111111111001010101100110011111010;
filter5[1][588] = 35'b00000000011011101010110011110001100;
filter5[1][589] = 35'b11111111101000110100111110101000000;
filter5[1][590] = 35'b11111110100000111110110010100010000;
filter5[1][591] = 35'b00000100110001110101010010100000000;
filter5[1][592] = 35'b00000100001111110000001001111000000;
filter5[1][593] = 35'b11111111111000100111111000001111010;
filter5[1][594] = 35'b11111111011000000110010100111010000;
filter5[1][595] = 35'b11111101011010010000111001100000000;
filter5[1][596] = 35'b11111110001011000110011100010000000;
filter5[1][597] = 35'b00000000011000011110010001111100000;
filter5[1][598] = 35'b00000000010100110000111100101100100;
filter5[1][599] = 35'b11111111010000101111101000110010000;
filter5[1][600] = 35'b00000011111001100010011001011100000;
filter5[1][601] = 35'b11111111101101000000010110111011100;
filter5[1][602] = 35'b00000000010111101011000100110001000;
filter5[1][603] = 35'b00000010101110101110100100110100000;
filter5[1][604] = 35'b00000010111100001110000100010000000;
filter5[1][605] = 35'b00000010001100000101000101110100000;
filter5[1][606] = 35'b11111000110010011101010100110000000;
filter5[1][607] = 35'b00000110101101101010111110101000000;
filter5[1][608] = 35'b00001000100100000110010000000000000;
filter5[1][609] = 35'b11111101101000000001110010111100000;
filter5[1][610] = 35'b00000011010111001010110101010100000;
filter5[1][611] = 35'b11111010111010011010000010101000000;
filter5[1][612] = 35'b00000001011001100101110101101000000;
filter5[1][613] = 35'b11111110100100100001100101001100000;
filter5[1][614] = 35'b11111110110001000000001000110000000;
filter5[1][615] = 35'b00000001010000011001110001100110000;
filter5[1][616] = 35'b00000011110100000011010010100000000;
filter5[1][617] = 35'b00000000100100110110001101010110000;
filter5[1][618] = 35'b11111111001001101100000100000110000;
filter5[1][619] = 35'b00000001011100001101000001000110000;
filter5[1][620] = 35'b11111110011110101011010000100100000;
filter5[1][621] = 35'b11111111110111111100001010111000000;
filter5[1][622] = 35'b11111110111100011011000100101100000;
filter5[1][623] = 35'b11111111011111101111111111000110000;
filter5[1][624] = 35'b11111110111011101010111000010100000;
filter5[1][625] = 35'b11111100000010111010001100010100000;
filter5[1][626] = 35'b00000000100001010011010110011110000;
filter5[1][627] = 35'b11111100000011100101101101110100000;
filter5[1][628] = 35'b11111101010110100100101110000100000;
filter5[1][629] = 35'b11111110000011110000011101000010000;
filter5[1][630] = 35'b00000000000111000100100001101001110;
filter5[1][631] = 35'b00000000101010100000111101111110000;
filter5[1][632] = 35'b00000000111110010000010111001000000;
filter5[1][633] = 35'b00000001000100001001111111110010000;
filter5[1][634] = 35'b00000000111011110011010100011110000;
filter5[1][635] = 35'b11111110010010100010100111010100000;
filter5[1][636] = 35'b11111101010000110000110000011000000;
filter5[1][637] = 35'b00000111010000010101110000100000000;
filter5[1][638] = 35'b00000010101111000001110010011000000;
filter5[1][639] = 35'b00000000011010011010000000111100100;
filter5[1][640] = 35'b00000101001100001001001111000000000;
filter5[1][641] = 35'b11111101010011100000111000011100000;
filter5[1][642] = 35'b11111110001100110100100111110000000;
filter5[1][643] = 35'b00000010011000111111110100011000000;
filter5[1][644] = 35'b11111111111100101001010011111010111;
filter5[1][645] = 35'b00000000011011101101010000110001000;
filter5[1][646] = 35'b11111110000011000101101001000100000;
filter5[1][647] = 35'b00000001000010000100000100001110000;
filter5[1][648] = 35'b11111100101110111010101100000000000;
filter5[1][649] = 35'b11111101110000010000000110001000000;
filter5[1][650] = 35'b11111110111011011010100000101110000;
filter5[1][651] = 35'b00000000110001100100100111110100000;
filter5[1][652] = 35'b00000000001111001000100101100001110;
filter5[1][653] = 35'b00000000101000010011101100010010000;
filter5[1][654] = 35'b11111111011011100011001000111011000;
filter5[1][655] = 35'b00000000010010010100001000001001100;
filter5[1][656] = 35'b11111001110101111011010001101000000;
filter5[1][657] = 35'b11111000100111001011110111101000000;
filter5[1][658] = 35'b11111000111110110011111111000000000;
filter5[1][659] = 35'b11111111001100010000101100000100000;
filter5[1][660] = 35'b11111101110000100101100110100000000;
filter5[1][661] = 35'b11111110001010010011110000100010000;
filter5[1][662] = 35'b11111100010000001100000100011000000;
filter5[1][663] = 35'b00000011011000110010011100010100000;
filter5[1][664] = 35'b00000100101010011111001111000000000;
filter5[1][665] = 35'b00000111111001001011010011111000000;
filter5[1][666] = 35'b11111110001110101110100000000100000;
filter5[1][667] = 35'b11111110010101001011000011011100000;
filter5[1][668] = 35'b11111110101010011110110011001110000;
filter5[1][669] = 35'b11111110111111001101110001100110000;
filter5[1][670] = 35'b00000001110111111010101011110100000;
filter5[1][671] = 35'b00000010111011001011011110001000000;
filter5[1][672] = 35'b00001010001111011111000001000000000;
filter5[1][673] = 35'b00000100100011011000100111111000000;
filter5[1][674] = 35'b00001001000011000100101110110000000;
filter5[1][675] = 35'b11111101101100111000011000101100000;
filter5[1][676] = 35'b00000011100010001100100000011000000;
filter5[1][677] = 35'b00000010100110011110000001111000000;
filter5[1][678] = 35'b11111110011101000001000000010100000;
filter5[1][679] = 35'b11111101010001010100110101111100000;
filter5[1][680] = 35'b11111110011001000111100101000100000;
filter5[1][681] = 35'b00000110011000000110000000000000000;
filter5[1][682] = 35'b00000101010011010110001010100000000;
filter5[1][683] = 35'b00000001000001100111011000000110000;
filter5[1][684] = 35'b11111111101100010000000001010000000;
filter5[1][685] = 35'b11111110101110011010000000101000000;
filter5[1][686] = 35'b11111101010111101011100111101000000;
filter5[1][687] = 35'b11111101010010011000001010111100000;
filter5[1][688] = 35'b11111011111010011000000010100000000;
filter5[1][689] = 35'b00000000000001010111101010111100111;
filter5[1][690] = 35'b11111101101111110101001100010100000;
filter5[1][691] = 35'b11111101101101111101011011101100000;
filter5[1][692] = 35'b00000000011000101110000011000000100;
filter5[1][693] = 35'b11111111010011100100010100100100000;
filter5[1][694] = 35'b11111110001000110101100010110010000;
filter5[1][695] = 35'b11111101111000000010110010011100000;
filter5[1][696] = 35'b11111100101110111101101111000000000;
filter5[1][697] = 35'b00000001101100111000100010010100000;
filter5[1][698] = 35'b00000010001000101001011110111000000;
filter5[1][699] = 35'b11111111001111010011111111110011000;
filter5[1][700] = 35'b11111111011011111111000101001001000;
filter5[1][701] = 35'b00000001001110010101000110000110000;
filter5[1][702] = 35'b11111111101111100010001111100100100;
filter5[1][703] = 35'b11111111001110001001011000100101000;
filter5[1][704] = 35'b11111101011101100101000010101000000;
filter5[1][705] = 35'b11111111000001111110110101000110000;
filter5[1][706] = 35'b00000001000010010111000011000000000;
filter5[1][707] = 35'b11111111111101111101110011011110111;
filter5[1][708] = 35'b11111111111101100101001010110111011;
filter5[1][709] = 35'b00000000101101010111010011010100000;
filter5[1][710] = 35'b00000001000011010000010111111110000;
filter5[1][711] = 35'b00000000010110100000100010100110000;
filter5[1][712] = 35'b00000000000100100001001010011110001;
filter5[1][713] = 35'b00000001111111010100101101110000000;
filter5[1][714] = 35'b00000100111001010110001100100000000;
filter5[1][715] = 35'b11111111010000011110010010011111000;
filter5[1][716] = 35'b11111101001111000000011100011100000;
filter5[1][717] = 35'b11111111111010101101101000111000100;
filter5[1][718] = 35'b00000001010000110011110110100100000;
filter5[1][719] = 35'b00000000011100000010111101000110100;
filter5[1][720] = 35'b11111111110111011010111000000100100;
filter5[1][721] = 35'b00000011010000101011100001100000000;
filter5[1][722] = 35'b00000000000000000001011000001100100;
filter5[1][723] = 35'b11111110000111001111001101110000000;
filter5[1][724] = 35'b00000001010010001001100101101110000;
filter5[1][725] = 35'b11111101001111101010010010011000000;
filter5[1][726] = 35'b11111111111111010111101100101101110;
filter5[1][727] = 35'b00000001000101000011011010111010000;
filter5[1][728] = 35'b00000001000011000101110000100000000;
filter5[1][729] = 35'b00000001110001000011010011100100000;
filter5[1][730] = 35'b00000100110010010100110011100000000;
filter5[1][731] = 35'b11111111101001110001100111110100000;
filter5[1][732] = 35'b11111101011000110001011000001100000;
filter5[1][733] = 35'b11111101110111010111100000000000000;
filter5[1][734] = 35'b11111100011101100111100111011100000;
filter5[1][735] = 35'b00000000011010110011011101111000100;
filter5[1][736] = 35'b11111101111001001010000001101100000;
filter5[1][737] = 35'b00000011001010001110111111110000000;
filter5[1][738] = 35'b00000110011010111001001000110000000;
filter5[1][739] = 35'b11111111111000101000010001010001101;
filter5[1][740] = 35'b00000000110000101101111100110001000;
filter5[1][741] = 35'b00000000101001100010001001010010000;
filter5[1][742] = 35'b11111001011110101001110101110000000;
filter5[1][743] = 35'b00000001100111101110011010101110000;
filter5[1][744] = 35'b11111100101111101010110011010000000;
filter5[1][745] = 35'b00000000001011101010100111001001110;
filter5[1][746] = 35'b00000100110000110011000011011000000;
filter5[1][747] = 35'b11111101000011000111110110011100000;
filter5[1][748] = 35'b11111101000100100111011011000000000;
filter5[1][749] = 35'b00000000101000111001101111011100000;
filter5[1][750] = 35'b11111110101001101011100001100100000;
filter5[1][751] = 35'b11111100000111001111100011111100000;
filter5[1][752] = 35'b11111010100011100010110010000000000;
filter5[1][753] = 35'b11111001101100010010101011000000000;
filter5[1][754] = 35'b11111101001010011100101001111100000;
filter5[1][755] = 35'b11111110001010100000110001100000000;
filter5[1][756] = 35'b11111111110010010100111111001111100;
filter5[1][757] = 35'b00000000110001111010101011100101000;
filter5[1][758] = 35'b11111101111110111000101010001100000;
filter5[1][759] = 35'b11111111001101101011110100011110000;
filter5[1][760] = 35'b11111110110001010010111011001010000;
filter5[1][761] = 35'b11111010010101011000001100000000000;
filter5[1][762] = 35'b00000010011010011011111100001000000;
filter5[1][763] = 35'b11111101101111110011100111110100000;
filter5[1][764] = 35'b00000010000110010000101111001000000;
filter5[1][765] = 35'b00000000111010010010000110111011000;
filter5[1][766] = 35'b11111101100111110101010101000000000;
filter5[1][767] = 35'b11111110101111011010011001001100000;
filter5[1][768] = 35'b00000100010000000001110100011000000;
filter5[1][769] = 35'b00000010011011010101101111100000000;
filter5[1][770] = 35'b00000000100100100000110110011111000;
filter5[1][771] = 35'b11111111101011101111000001010101000;
filter5[1][772] = 35'b11111111111011001100000110000010111;
filter5[1][773] = 35'b00000001010110000000111001111000000;
filter5[1][774] = 35'b11111101111001001011011010011100000;
filter5[1][775] = 35'b00000010010001001011000110001100000;
filter5[1][776] = 35'b00000100001000101100010000010000000;
filter5[1][777] = 35'b00000000111000101000101011000010000;
filter5[1][778] = 35'b11111001111110001110101001011000000;
filter5[1][779] = 35'b00000100100010001100010111101000000;
filter5[1][780] = 35'b11111111000010111110110000110000000;
filter5[1][781] = 35'b11111111001001011101111011011001000;
filter5[1][782] = 35'b00000000001001001101000011111100000;
filter5[1][783] = 35'b00000000100100010111000101100101000;
filter5[1][784] = 35'b00000000111011110110111010101000000;
filter5[1][785] = 35'b00000001000101001100011100010000000;
filter5[1][786] = 35'b11110111110110110001111110100000000;
filter5[1][787] = 35'b00000010010100011011101100011100000;
filter5[1][788] = 35'b00000010011101001111110011000100000;
filter5[1][789] = 35'b11111010101101011111010101100000000;
filter5[1][790] = 35'b00000011001100101100110000010000000;
filter5[1][791] = 35'b00000000101000000011001101101110000;
filter5[1][792] = 35'b11111111101001100000110100101001000;
filter5[1][793] = 35'b11111111011110000101010100010000000;
filter5[1][794] = 35'b11111101010110111011001011000100000;
filter5[1][795] = 35'b11111110001101001111110110111000000;
filter5[1][796] = 35'b00000011010001101101100100111100000;
filter5[1][797] = 35'b11111111101110010111100101110110100;
filter5[1][798] = 35'b00000110001100011110101110111000000;
filter5[1][799] = 35'b11111011001001001011000010100000000;
filter5[1][800] = 35'b00000100010011011011000000001000000;
filter5[1][801] = 35'b00001000110000111100111001000000000;
filter5[1][802] = 35'b00000001010100101100011010011110000;
filter5[1][803] = 35'b00000101011101100100100010000000000;
filter5[1][804] = 35'b11111101011011000110100111111000000;
filter5[1][805] = 35'b11111110101001011111110111011110000;
filter5[1][806] = 35'b00000001101101000111011111000110000;
filter5[1][807] = 35'b11111011100011000000100001010000000;
filter5[1][808] = 35'b00000010001110010111100110000000000;
filter5[1][809] = 35'b00000100001111101001101010100000000;
filter5[1][810] = 35'b00000010110100011001100100010100000;
filter5[1][811] = 35'b00000010100011011101010110111000000;
filter5[1][812] = 35'b00000001111110101010010101000100000;
filter5[1][813] = 35'b11111110100011100010111110001000000;
filter5[1][814] = 35'b00000001010100100010100010011010000;
filter5[1][815] = 35'b11111101010000010110000111110100000;
filter5[1][816] = 35'b11111111101011010000001111011001100;
filter5[1][817] = 35'b11111101000110101100001010100000000;
filter5[1][818] = 35'b11111101111000111110111010111000000;
filter5[1][819] = 35'b00000000001000100110110001001001100;
filter5[1][820] = 35'b11111100011011001001111001011100000;
filter5[1][821] = 35'b11111100011100011111100010110000000;
filter5[1][822] = 35'b11111101010101010001101000011100000;
filter5[1][823] = 35'b00000000111010100001111010011000000;
filter5[1][824] = 35'b11111011100100011111110110000000000;
filter5[1][825] = 35'b00000101110110010111001000100000000;
filter5[1][826] = 35'b00000001110101111100111110011100000;
filter5[1][827] = 35'b11111110101111001100000010001100000;
filter5[1][828] = 35'b11111011111110101000001001110000000;
filter5[1][829] = 35'b11111100110100011011011001001000000;
filter5[1][830] = 35'b11111111100101001011100001000000100;
filter5[1][831] = 35'b11111101100110000000000010000000000;
filter5[1][832] = 35'b00000000010111110111111000110101000;
filter5[1][833] = 35'b11111110001000000010100000101110000;
filter5[1][834] = 35'b11111111000111111001110110010000000;
filter5[1][835] = 35'b11111110111001101110010111011010000;
filter5[1][836] = 35'b11111111010001011111010011010011000;
filter5[1][837] = 35'b00000001100110001110011011000000000;
filter5[1][838] = 35'b00000000001011010100111111000101010;
filter5[1][839] = 35'b00000000000100011011000001110010100;
filter5[1][840] = 35'b11111110111100000010010010000100000;
filter5[1][841] = 35'b11111110111101001100100111101010000;
filter5[1][842] = 35'b00000000110111110100011110111100000;
filter5[1][843] = 35'b11111110011000110100010110100010000;
filter5[1][844] = 35'b11111111110101110011010000100110000;
filter5[1][845] = 35'b11111111101010100010111111110010000;
filter5[1][846] = 35'b11111111110111011111111000101011010;
filter5[1][847] = 35'b11111111100100111101101101110111100;
filter5[1][848] = 35'b00000010000000111111101100100100000;
filter5[1][849] = 35'b00000100000010100010110110110000000;
filter5[1][850] = 35'b00000000000100001100011011011000011;
filter5[1][851] = 35'b11111101000100000000011010100000000;
filter5[1][852] = 35'b00000010100010010110110111100000000;
filter5[1][853] = 35'b11111010100001001110100111111000000;
filter5[1][854] = 35'b00000001101101000000111010000010000;
filter5[1][855] = 35'b00000000010010011001001011000110000;
filter5[1][856] = 35'b11111100110101011010000101000100000;
filter5[1][857] = 35'b00000000110101111101000010101001000;
filter5[1][858] = 35'b00000010000101001011011001010000000;
filter5[1][859] = 35'b00000000011110000010001100111110000;
filter5[1][860] = 35'b00000000101010010011001001111110000;
filter5[1][861] = 35'b11111010001111001000101100100000000;
filter5[1][862] = 35'b11111101101000111001001111000100000;
filter5[1][863] = 35'b00000001110001100101100001111110000;
filter5[1][864] = 35'b11111110100111000000100000111110000;
filter5[1][865] = 35'b00000010001101001100101100110100000;
filter5[1][866] = 35'b00000100111100011011100110110000000;
filter5[1][867] = 35'b11111101011001101101111101011100000;
filter5[1][868] = 35'b00000010100001101010011001111000000;
filter5[1][869] = 35'b11110101101011101111001111000000000;
filter5[1][870] = 35'b00000001111010101001101110111010000;
filter5[1][871] = 35'b00000001110110101101001100011100000;
filter5[1][872] = 35'b11111110001100111101111101001100000;
filter5[1][873] = 35'b11111111111010010100111101011101001;
filter5[1][874] = 35'b00000010111011100110011101010000000;
filter5[1][875] = 35'b11111011100100000011001000001000000;
filter5[1][876] = 35'b11111111001011001000111010001111000;
filter5[1][877] = 35'b00000010010111110010011100001100000;
filter5[1][878] = 35'b11111000001100010010100101001000000;
filter5[1][879] = 35'b00000000011111010101111110101111000;
filter5[1][880] = 35'b11111101000101110011000011111100000;
filter5[1][881] = 35'b11111101111000111000101111100000000;
filter5[1][882] = 35'b00000000000110011111011111100000011;
filter5[1][883] = 35'b11111111100011110000101100011110100;
filter5[1][884] = 35'b11111011011000011111010011100000000;
filter5[1][885] = 35'b11111101010001100001000010111000000;
filter5[1][886] = 35'b11111101000000011001111001111100000;
filter5[1][887] = 35'b11111111110101111101110001010001010;
filter5[1][888] = 35'b11111100010000101011001111101100000;
filter5[1][889] = 35'b11111111111011100101011001001010101;
filter5[1][890] = 35'b11111111101011000100010011101101100;
filter5[1][891] = 35'b11111100111000101111110010110100000;
filter5[1][892] = 35'b00000011111100000001100100101100000;
filter5[1][893] = 35'b00000100000000100011100100011000000;
filter5[1][894] = 35'b11111101000110100110010000110000000;
filter5[1][895] = 35'b11111101111101001000111011100100000;
filter5[1][896] = 35'b11111010100000111110110011101000000;
filter5[1][897] = 35'b11111000100011110000001101100000000;
filter5[1][898] = 35'b11110011000101101100110011100000000;
filter5[1][899] = 35'b11111100011010001010101000101100000;
filter5[1][900] = 35'b11111111111011010001111110011010001;
filter5[1][901] = 35'b00000000000011111000001111100111110;
filter5[1][902] = 35'b11111101111111101001110100001100000;
filter5[1][903] = 35'b00000101011001101101100010111000000;
filter5[1][904] = 35'b11111010001100111001110010010000000;
filter5[1][905] = 35'b00000001010001011101000001000000000;
filter5[1][906] = 35'b00000101011000011110001001110000000;
filter5[1][907] = 35'b11111011010001101010001001110000000;
filter5[1][908] = 35'b11110001011100010110101010010000000;
filter5[1][909] = 35'b11111101100101100101101010011100000;
filter5[1][910] = 35'b11111011010101110101010101011000000;
filter5[1][911] = 35'b11111110011101110100011000101000000;
filter5[1][912] = 35'b00000000100011110001000111110111000;
filter5[1][913] = 35'b00000000010011101110110001010010100;
filter5[1][914] = 35'b00000001101101001110000101110110000;
filter5[1][915] = 35'b00000000010000100100100001010100000;
filter5[1][916] = 35'b00000001001000011001010110010010000;
filter5[1][917] = 35'b11110010000100010010011001010000000;
filter5[1][918] = 35'b11111010100101000101011110100000000;
filter5[1][919] = 35'b11111101000011001000100101101100000;
filter5[1][920] = 35'b00000010110110010011000000011100000;
filter5[1][921] = 35'b00000010000011000110101101001000000;
filter5[1][922] = 35'b00000011000011010011101000111000000;
filter5[1][923] = 35'b11111110100001011011011001101010000;
filter5[1][924] = 35'b00000000110100000111000111001100000;
filter5[1][925] = 35'b11111000000010001101101110011000000;
filter5[1][926] = 35'b11111011110110001101010101110000000;
filter5[1][927] = 35'b11111111010011001110111001111011000;
filter5[1][928] = 35'b11111101111001000001100100110000000;
filter5[1][929] = 35'b00000011110100010011101110110100000;
filter5[1][930] = 35'b00000010010001101000010011001100000;
filter5[1][931] = 35'b11111111110110111001001101100111010;
filter5[1][932] = 35'b00000001001110100100000100101100000;
filter5[1][933] = 35'b11110110110010110110100011000000000;
filter5[1][934] = 35'b11110111110100100011101110100000000;
filter5[1][935] = 35'b11111001100110001011110001110000000;
filter5[1][936] = 35'b11111110011110110000011100011100000;
filter5[1][937] = 35'b11111001111011000000010001010000000;
filter5[1][938] = 35'b11111111111100100011000110111000110;
filter5[1][939] = 35'b11111010010011101000111011011000000;
filter5[1][940] = 35'b11111110101110000110100101011110000;
filter5[1][941] = 35'b00000100000000101101110111110000000;
filter5[1][942] = 35'b11110111010011000100101011100000000;
filter5[1][943] = 35'b00000000000110101110110010011101100;
filter5[1][944] = 35'b11110011111011101000011010110000000;
filter5[1][945] = 35'b00000010111000001110011011111000000;
filter5[1][946] = 35'b00000011110100000110000001100000000;
filter5[1][947] = 35'b00000000111101001100111110011011000;
filter5[1][948] = 35'b11111011110111001100110110000000000;
filter5[1][949] = 35'b00000001111001100010100100101110000;
filter5[1][950] = 35'b11101100010010011010010110100000000;
filter5[1][951] = 35'b11111111001101001000011001111111000;
filter5[1][952] = 35'b11111000100010000110010001010000000;
filter5[1][953] = 35'b11111001111011011010001100111000000;
filter5[1][954] = 35'b11111100100001101111100110111100000;
filter5[1][955] = 35'b11111010011011011010000010010000000;
filter5[1][956] = 35'b00000001011110110100000000000110000;
filter5[1][957] = 35'b00000000010001100111111000001010000;
filter5[1][958] = 35'b11110100000101001010011000100000000;
filter5[1][959] = 35'b11111000111110001100010000000000000;
filter5[1][960] = 35'b00001000010110011000011010100000000;
filter5[1][961] = 35'b11111110000111011010011000011010000;
filter5[1][962] = 35'b11111010001001101111101110100000000;
filter5[1][963] = 35'b11111010000001110100111000111000000;
filter5[1][964] = 35'b11111100011011101110000110001000000;
filter5[1][965] = 35'b00000001001000110001001110111000000;
filter5[1][966] = 35'b00000110001100000110100111101000000;
filter5[1][967] = 35'b11111111011100011100110111101111000;
filter5[1][968] = 35'b11111101110011101010010100001000000;
filter5[1][969] = 35'b00000010001010001000011010000000000;
filter5[1][970] = 35'b00000110101001010000111110101000000;
filter5[1][971] = 35'b00000011011001011001010001110000000;
filter5[1][972] = 35'b11111011011111110101111100011000000;
filter5[1][973] = 35'b11111000001101101001101101010000000;
filter5[1][974] = 35'b00000001011010101011110011101000000;
filter5[1][975] = 35'b00000010010011000111101101001100000;
filter5[1][976] = 35'b00000011000001110101110010101000000;
filter5[1][977] = 35'b00000001011000100110000101001110000;
filter5[1][978] = 35'b00000001011111001011100100000000000;
filter5[1][979] = 35'b00000010001010001110111000010000000;
filter5[1][980] = 35'b00000011100001111111000110010100000;
filter5[1][981] = 35'b11111110100001100101100010001000000;
filter5[1][982] = 35'b11110111011111000111010100110000000;
filter5[1][983] = 35'b11111101001110011001010010001100000;
filter5[1][984] = 35'b00000000010011001010001001100111000;
filter5[1][985] = 35'b11111111110111001111000100111010000;
filter5[1][986] = 35'b00000000101101011110001110101111000;
filter5[1][987] = 35'b00000011001000011100110000001000000;
filter5[1][988] = 35'b11111100111100010010011010110000000;
filter5[1][989] = 35'b11111100001110110101100001011100000;
filter5[1][990] = 35'b11111001011100011101001110111000000;
filter5[1][991] = 35'b00000000010001001100110010110111000;
filter5[1][992] = 35'b00000110010100110010101001101000000;
filter5[1][993] = 35'b00000011101000011101001011010000000;
filter5[1][994] = 35'b11111100001100010011000011111100000;
filter5[1][995] = 35'b00000000110011010111100110000111000;
filter5[1][996] = 35'b00000011010110101111101101100000000;
filter5[1][997] = 35'b00000101000000000010010111100000000;
filter5[1][998] = 35'b00000001010001110111010000101110000;
filter5[1][999] = 35'b11111101000110100100001101001000000;
filter5[1][1000] = 35'b00001000100010101110100011110000000;
filter5[1][1001] = 35'b00000110010111010011111101000000000;
filter5[1][1002] = 35'b11111011110011111001110101111000000;
filter5[1][1003] = 35'b00000000110101111101100001101111000;
filter5[1][1004] = 35'b11110010100101101100100101000000000;
filter5[1][1005] = 35'b11111100111110011001110100010100000;
filter5[1][1006] = 35'b11111101101101110001111001110100000;
filter5[1][1007] = 35'b00000010111010001110110001011100000;
filter5[1][1008] = 35'b00000001010000000000001100010010000;
filter5[1][1009] = 35'b11110110110100000111011100010000000;
filter5[1][1010] = 35'b11100111100001001100001000000000000;
filter5[1][1011] = 35'b11110001000100011011111000000000000;
filter5[1][1012] = 35'b11111011101111100000001010011000000;
filter5[1][1013] = 35'b00000001101001010111000110010010000;
filter5[1][1014] = 35'b00000010101010010110111110010000000;
filter5[1][1015] = 35'b11111011110010101001100100100000000;
filter5[1][1016] = 35'b11111100100010010100010101101000000;
filter5[1][1017] = 35'b11111111100001000111111100001001100;
filter5[1][1018] = 35'b11111100101100001001100100101000000;
filter5[1][1019] = 35'b11111011000110000001000101100000000;
filter5[1][1020] = 35'b00000010111001110110110111000000000;
filter5[1][1021] = 35'b11111101011101010111011001010100000;
filter5[1][1022] = 35'b11111011010111110101101110001000000;
filter5[1][1023] = 35'b11111011101110110101010110110000000;
filter5[2][0] = 35'b00000000000011100100010001101011100;
filter5[2][1] = 35'b11111001010000110010010010010000000;
filter5[2][2] = 35'b11111100011010011110100001110100000;
filter5[2][3] = 35'b11111101000100100010111001011000000;
filter5[2][4] = 35'b11111100010100000011101111110100000;
filter5[2][5] = 35'b11111110001001000111101100000000000;
filter5[2][6] = 35'b00000000011011000001010100100111100;
filter5[2][7] = 35'b00000000000110110101110111001010101;
filter5[2][8] = 35'b00000111001110001111111111000000000;
filter5[2][9] = 35'b00000010000011010010100011101000000;
filter5[2][10] = 35'b11111101101100110101001011101000000;
filter5[2][11] = 35'b11111000100010100111011001001000000;
filter5[2][12] = 35'b00000011001001011010001000000000000;
filter5[2][13] = 35'b11111011000011100000100100111000000;
filter5[2][14] = 35'b00000001000001001111000111110000000;
filter5[2][15] = 35'b00000100011111111100000101000000000;
filter5[2][16] = 35'b00000010000100011011101010011000000;
filter5[2][17] = 35'b00000011111010110100110000000000000;
filter5[2][18] = 35'b11111100101001100110001101100100000;
filter5[2][19] = 35'b00000001000111010101101011110110000;
filter5[2][20] = 35'b11111111100010100010110101100010100;
filter5[2][21] = 35'b11111011010101100010000001110000000;
filter5[2][22] = 35'b00000011001111101111001110101100000;
filter5[2][23] = 35'b00000011110000000101101000111100000;
filter5[2][24] = 35'b00000011100000011100100101110100000;
filter5[2][25] = 35'b00000011111100011001110011010000000;
filter5[2][26] = 35'b00000011011111101000110100000100000;
filter5[2][27] = 35'b11111111010000010011110010100000000;
filter5[2][28] = 35'b11111111111111011110111010001110000;
filter5[2][29] = 35'b00000001101110111001000001101100000;
filter5[2][30] = 35'b11111011000001111110110110111000000;
filter5[2][31] = 35'b11111011101000000111000010100000000;
filter5[2][32] = 35'b00000000011101111000000101110101100;
filter5[2][33] = 35'b11111110100100011100000010011000000;
filter5[2][34] = 35'b11111111001001100111111000111011000;
filter5[2][35] = 35'b00000001001011010111111010000000000;
filter5[2][36] = 35'b00000011110111100111011001001000000;
filter5[2][37] = 35'b00000011111010001110110000010000000;
filter5[2][38] = 35'b00000101101010111011000101010000000;
filter5[2][39] = 35'b11111100100000011110101110010000000;
filter5[2][40] = 35'b00000001010011101101001001111100000;
filter5[2][41] = 35'b00000000010100111010100010111111000;
filter5[2][42] = 35'b11111111011100100001011101001110000;
filter5[2][43] = 35'b11111111111111000101010011011111110;
filter5[2][44] = 35'b11111010010100010110000001010000000;
filter5[2][45] = 35'b11111111011011111010110001110100000;
filter5[2][46] = 35'b00000110110110001000111000100000000;
filter5[2][47] = 35'b11111101111111001110111000100000000;
filter5[2][48] = 35'b11111100011010101011000001011100000;
filter5[2][49] = 35'b11111110001001000010010111100000000;
filter5[2][50] = 35'b11111111000011110101000101110000000;
filter5[2][51] = 35'b11111111101111100100000010100011100;
filter5[2][52] = 35'b11111100011010010101011000100100000;
filter5[2][53] = 35'b00001000111000000010111111110000000;
filter5[2][54] = 35'b11111011110000011110010001000000000;
filter5[2][55] = 35'b11111110001111011011010001110110000;
filter5[2][56] = 35'b11111100111000101011101001111100000;
filter5[2][57] = 35'b00000101001100000101011100010000000;
filter5[2][58] = 35'b00000011111011111100001000011000000;
filter5[2][59] = 35'b11111101110001111101111010010000000;
filter5[2][60] = 35'b11111111000110110011010111011011000;
filter5[2][61] = 35'b11111010000000011010100000001000000;
filter5[2][62] = 35'b00000010110110011000011100110000000;
filter5[2][63] = 35'b11111110101000111110111010111000000;
filter5[2][64] = 35'b11111110000100101101000001111010000;
filter5[2][65] = 35'b11111101011110100001110001100000000;
filter5[2][66] = 35'b11111110111011010101110001100110000;
filter5[2][67] = 35'b11111010111000000001001010111000000;
filter5[2][68] = 35'b11111101101101001010011011100100000;
filter5[2][69] = 35'b11111101000000111000001001110100000;
filter5[2][70] = 35'b11111111000101011010100101010000000;
filter5[2][71] = 35'b11111110111011000010101110100000000;
filter5[2][72] = 35'b00000000110111001001101001100011000;
filter5[2][73] = 35'b00000001010001101010010000000000000;
filter5[2][74] = 35'b00000001110010100011000011011100000;
filter5[2][75] = 35'b11111110010101000000001000000010000;
filter5[2][76] = 35'b00000010001100111010101001111000000;
filter5[2][77] = 35'b00000000001100000001010000101101010;
filter5[2][78] = 35'b11111111000110001011001001101010000;
filter5[2][79] = 35'b11111110001010100000000001010010000;
filter5[2][80] = 35'b11111110100010100110110101101000000;
filter5[2][81] = 35'b00000010000001100110010111001000000;
filter5[2][82] = 35'b11111100100110110110111011010100000;
filter5[2][83] = 35'b11111111101000111110100101100101100;
filter5[2][84] = 35'b00000000011001101001101111011111000;
filter5[2][85] = 35'b11111100111101000100001101100000000;
filter5[2][86] = 35'b11111111001001101011011001110000000;
filter5[2][87] = 35'b00000000101010111010001101110001000;
filter5[2][88] = 35'b00000000110111010111101001100001000;
filter5[2][89] = 35'b00000010000110101000110101110100000;
filter5[2][90] = 35'b00000010001010111001011000101100000;
filter5[2][91] = 35'b11111110011111100111100100011110000;
filter5[2][92] = 35'b11111101011001000100000000111100000;
filter5[2][93] = 35'b00000001000000001011011100001000000;
filter5[2][94] = 35'b11111111011011110010110001101110000;
filter5[2][95] = 35'b11111111111001100111101111000110100;
filter5[2][96] = 35'b00000000100000111101000101000011000;
filter5[2][97] = 35'b11111100110110001011011100001000000;
filter5[2][98] = 35'b11111100010100000011011011001000000;
filter5[2][99] = 35'b00000010110000000101001010011000000;
filter5[2][100] = 35'b00000010111001001111111101111000000;
filter5[2][101] = 35'b00000100010010011000000110110000000;
filter5[2][102] = 35'b00000010010110011000001100111000000;
filter5[2][103] = 35'b00000010011010101100101110011100000;
filter5[2][104] = 35'b00000000010110010010111110101000000;
filter5[2][105] = 35'b00000000110000101011111011110110000;
filter5[2][106] = 35'b11111101000110010101001001101000000;
filter5[2][107] = 35'b11111110001011000110011111100100000;
filter5[2][108] = 35'b11111101100111100111000111011100000;
filter5[2][109] = 35'b00000010101011100110100001000000000;
filter5[2][110] = 35'b11111010010100110001011101001000000;
filter5[2][111] = 35'b11111101011101010000010100100100000;
filter5[2][112] = 35'b11111100111100000000010011110100000;
filter5[2][113] = 35'b11111111000010111001010100001110000;
filter5[2][114] = 35'b00000001010010010001111110001100000;
filter5[2][115] = 35'b11111111101101001011100101111010100;
filter5[2][116] = 35'b11111101011010111000110010010100000;
filter5[2][117] = 35'b00000010101101111001101001000100000;
filter5[2][118] = 35'b11111100110100010001110110101100000;
filter5[2][119] = 35'b00000000000010001001111001010111111;
filter5[2][120] = 35'b00000010110101100001101110011100000;
filter5[2][121] = 35'b00000110011111111010001111011000000;
filter5[2][122] = 35'b00000001101111110001100110001000000;
filter5[2][123] = 35'b11111100101011000001101001101100000;
filter5[2][124] = 35'b11111110110001101111100100001010000;
filter5[2][125] = 35'b11111111010100010000101000011011000;
filter5[2][126] = 35'b00000010011011110110110100110000000;
filter5[2][127] = 35'b11111101010001101100010001000100000;
filter5[2][128] = 35'b11111111001111111010111101010001000;
filter5[2][129] = 35'b11110101001100001001010110110000000;
filter5[2][130] = 35'b11110100010111010000100001010000000;
filter5[2][131] = 35'b11110011011101011011110000010000000;
filter5[2][132] = 35'b11110011101101011101001011100000000;
filter5[2][133] = 35'b11101101001011110110001010000000000;
filter5[2][134] = 35'b11101101110101111110110011100000000;
filter5[2][135] = 35'b11111000001010100000111101100000000;
filter5[2][136] = 35'b11111111011101001010111010010011000;
filter5[2][137] = 35'b11110010000110110001101111100000000;
filter5[2][138] = 35'b00000010011100010010000111100000000;
filter5[2][139] = 35'b11110011110110011101010110110000000;
filter5[2][140] = 35'b00000011001000101000011011100000000;
filter5[2][141] = 35'b11111101100100110111000000100100000;
filter5[2][142] = 35'b00000001101101001001100101010110000;
filter5[2][143] = 35'b00000011101011100000110011110100000;
filter5[2][144] = 35'b00000010111011100001101110011000000;
filter5[2][145] = 35'b00000101110110001100111111011000000;
filter5[2][146] = 35'b11111010101111101001110010000000000;
filter5[2][147] = 35'b11111111100101101101100011011110000;
filter5[2][148] = 35'b11111110100010000011100110100110000;
filter5[2][149] = 35'b11111110100001001000110001001110000;
filter5[2][150] = 35'b00000001100110110100101101010000000;
filter5[2][151] = 35'b00000010001011010010001000001000000;
filter5[2][152] = 35'b00000100011111000010110001110000000;
filter5[2][153] = 35'b00000000111001011011010010100000000;
filter5[2][154] = 35'b00000001110000101010111000100010000;
filter5[2][155] = 35'b00000010100101000011101000111000000;
filter5[2][156] = 35'b11111101010000110111101010010000000;
filter5[2][157] = 35'b00000101000100010110001001010000000;
filter5[2][158] = 35'b00000010000011111110000111101100000;
filter5[2][159] = 35'b00000001100010001101010100101110000;
filter5[2][160] = 35'b11110111011111011110100010110000000;
filter5[2][161] = 35'b11110001010110011001000011000000000;
filter5[2][162] = 35'b11111011011011101110010111100000000;
filter5[2][163] = 35'b11111110000101110111010011000110000;
filter5[2][164] = 35'b00000000110101110010000101111000000;
filter5[2][165] = 35'b00001000110110100000001001110000000;
filter5[2][166] = 35'b00000000101000000000001000010001000;
filter5[2][167] = 35'b00001000011100111101100011110000000;
filter5[2][168] = 35'b00001000100000000101000111110000000;
filter5[2][169] = 35'b11111111001011101010010100010110000;
filter5[2][170] = 35'b11111101100110000010111110011100000;
filter5[2][171] = 35'b11110100001101100110110101000000000;
filter5[2][172] = 35'b11111000101110001110111111000000000;
filter5[2][173] = 35'b00000001001110011100011110110110000;
filter5[2][174] = 35'b11110111010100000100001110100000000;
filter5[2][175] = 35'b00001001111101011000010101000000000;
filter5[2][176] = 35'b00000101000000011100100011110000000;
filter5[2][177] = 35'b11111100010110001010011111001100000;
filter5[2][178] = 35'b11111001101101101010110110110000000;
filter5[2][179] = 35'b11111010000000000000000000101000000;
filter5[2][180] = 35'b11110000011111110000100111100000000;
filter5[2][181] = 35'b11110111000100000010010111100000000;
filter5[2][182] = 35'b11111010100110001001100100011000000;
filter5[2][183] = 35'b11111001101000000100001001101000000;
filter5[2][184] = 35'b11111101010011000111010010111100000;
filter5[2][185] = 35'b00000001101100111001110010010110000;
filter5[2][186] = 35'b11111100000111001100101001000100000;
filter5[2][187] = 35'b11111101100101101100101101010000000;
filter5[2][188] = 35'b11111100110100000111000010101100000;
filter5[2][189] = 35'b11111101100001001011011111010000000;
filter5[2][190] = 35'b11111001101001110111010011111000000;
filter5[2][191] = 35'b11110110010111100100110100110000000;
filter5[2][192] = 35'b11111010011000101100001011000000000;
filter5[2][193] = 35'b11110011111011001000101010100000000;
filter5[2][194] = 35'b00000010110010010100100010110000000;
filter5[2][195] = 35'b11111010010100010110001101101000000;
filter5[2][196] = 35'b11111001101100100001101100101000000;
filter5[2][197] = 35'b11110011011001110111011111010000000;
filter5[2][198] = 35'b11111001010010011101010110011000000;
filter5[2][199] = 35'b11111000010001011110101011010000000;
filter5[2][200] = 35'b00001000110011000000100110100000000;
filter5[2][201] = 35'b11111011101110101001010001001000000;
filter5[2][202] = 35'b11111110000111011101101000011010000;
filter5[2][203] = 35'b00000000111111100111011111101000000;
filter5[2][204] = 35'b11110110001100111101111111000000000;
filter5[2][205] = 35'b11111110001011110000101101001000000;
filter5[2][206] = 35'b00000000110111011011011000000101000;
filter5[2][207] = 35'b00000000000101110101010101101110000;
filter5[2][208] = 35'b00000011100111010111001110110000000;
filter5[2][209] = 35'b11111000110011000100100100111000000;
filter5[2][210] = 35'b11110111001000101111100101000000000;
filter5[2][211] = 35'b11111101100001001100000000011000000;
filter5[2][212] = 35'b00000010000001111100101100111000000;
filter5[2][213] = 35'b11110111011110111000101111110000000;
filter5[2][214] = 35'b11111100011110111011001001001100000;
filter5[2][215] = 35'b11111111110101100111011111000000110;
filter5[2][216] = 35'b00000100100011000010111110110000000;
filter5[2][217] = 35'b11111100110011110111101000010100000;
filter5[2][218] = 35'b11110100010100011011001010110000000;
filter5[2][219] = 35'b00000100110010100100100010101000000;
filter5[2][220] = 35'b11111110000000011100110001101100000;
filter5[2][221] = 35'b00000000010011000011111100001110100;
filter5[2][222] = 35'b00000011010011100100000011011100000;
filter5[2][223] = 35'b00000001010001111110101011100110000;
filter5[2][224] = 35'b11111001001001101111010100010000000;
filter5[2][225] = 35'b00000010010100110111101000101000000;
filter5[2][226] = 35'b11111101111000100010011100011100000;
filter5[2][227] = 35'b00000001100101111010101010111100000;
filter5[2][228] = 35'b00000010000111101011011111001100000;
filter5[2][229] = 35'b00000001011001101011011011010100000;
filter5[2][230] = 35'b11111111100111001010001001011101100;
filter5[2][231] = 35'b11111100101111100101010111100100000;
filter5[2][232] = 35'b11111000110011111111011101111000000;
filter5[2][233] = 35'b11111011100000110111010001101000000;
filter5[2][234] = 35'b11111110111100111110011101010010000;
filter5[2][235] = 35'b11111101001101010001101001000000000;
filter5[2][236] = 35'b11111011011011010110111100010000000;
filter5[2][237] = 35'b00000001000111011111001010010110000;
filter5[2][238] = 35'b00000100011101100100111110000000000;
filter5[2][239] = 35'b00000000110000011000000000000000000;
filter5[2][240] = 35'b11110010100111011010100101110000000;
filter5[2][241] = 35'b11111110000011110100101111000100000;
filter5[2][242] = 35'b11111111001011011010111111011111000;
filter5[2][243] = 35'b00000010010011001010000101110000000;
filter5[2][244] = 35'b11111101100110010010000111010000000;
filter5[2][245] = 35'b11111100011100100110010001101100000;
filter5[2][246] = 35'b11111101111000010001010010100100000;
filter5[2][247] = 35'b11111100111001000000110000001000000;
filter5[2][248] = 35'b11110111110001111010011110010000000;
filter5[2][249] = 35'b00001100000010010111101101110000000;
filter5[2][250] = 35'b00000010100100000110101111110000000;
filter5[2][251] = 35'b11111111111011110101101011001000000;
filter5[2][252] = 35'b11111011110010111100010110101000000;
filter5[2][253] = 35'b11111111100000011100111110000011100;
filter5[2][254] = 35'b11111110110111001010110101101010000;
filter5[2][255] = 35'b11111111011000100111110011110110000;
filter5[2][256] = 35'b11111110011010111011100101011010000;
filter5[2][257] = 35'b00000001110010010101101000011110000;
filter5[2][258] = 35'b11111110010100000111000011101100000;
filter5[2][259] = 35'b11111110101001010000101101110000000;
filter5[2][260] = 35'b11111011101101100100101011110000000;
filter5[2][261] = 35'b11111010100101101101111111010000000;
filter5[2][262] = 35'b11111100111111100001000100110100000;
filter5[2][263] = 35'b11111111000111111100100011011001000;
filter5[2][264] = 35'b00000000000101111101000011011111011;
filter5[2][265] = 35'b11111111011110011001011000110111000;
filter5[2][266] = 35'b11111110010000111001011011110110000;
filter5[2][267] = 35'b11111101111101010001100110111100000;
filter5[2][268] = 35'b11111110011011100110001011101010000;
filter5[2][269] = 35'b00000000010011101110000011101111000;
filter5[2][270] = 35'b11110110100111011011110001000000000;
filter5[2][271] = 35'b11110111101011011010010000100000000;
filter5[2][272] = 35'b11111010110100011100111000001000000;
filter5[2][273] = 35'b11111010110100111011001011110000000;
filter5[2][274] = 35'b11111000111010111010010011000000000;
filter5[2][275] = 35'b00000000100000100111110001001101000;
filter5[2][276] = 35'b11111101111101110110111011101000000;
filter5[2][277] = 35'b11111110010101100011000111100010000;
filter5[2][278] = 35'b00000000110001101011010010010000000;
filter5[2][279] = 35'b00001110000110101100101111000000000;
filter5[2][280] = 35'b11110111101110010010010001010000000;
filter5[2][281] = 35'b11110001000111101001000110110000000;
filter5[2][282] = 35'b11110110100110000000011010100000000;
filter5[2][283] = 35'b00000000000010110110111111110101001;
filter5[2][284] = 35'b00000010000111101110011111010100000;
filter5[2][285] = 35'b00000001000000110110111010110100000;
filter5[2][286] = 35'b00000110001111010010001110101000000;
filter5[2][287] = 35'b00000001000001001110001110011000000;
filter5[2][288] = 35'b11111101011011101000010101101100000;
filter5[2][289] = 35'b11111001111011100000101000110000000;
filter5[2][290] = 35'b11111011011000001000110100001000000;
filter5[2][291] = 35'b11111011110000110010000111111000000;
filter5[2][292] = 35'b00000000010111100100010100000001000;
filter5[2][293] = 35'b11111110101001100110010111001110000;
filter5[2][294] = 35'b00000001011111110110010111110010000;
filter5[2][295] = 35'b11111001010100011110100000001000000;
filter5[2][296] = 35'b11111011110000000000001011110000000;
filter5[2][297] = 35'b11110111101110101011111101010000000;
filter5[2][298] = 35'b00000001010000001101001110010110000;
filter5[2][299] = 35'b11111011001000100010011001011000000;
filter5[2][300] = 35'b11111111101011000000110011101110000;
filter5[2][301] = 35'b00000000000000001101001101100110100;
filter5[2][302] = 35'b11111101000001101111111101010100000;
filter5[2][303] = 35'b11111010011110100000110100101000000;
filter5[2][304] = 35'b11110101011001100101010100000000000;
filter5[2][305] = 35'b11111101101011001100010100111100000;
filter5[2][306] = 35'b11110101100011111000100110000000000;
filter5[2][307] = 35'b11110110101111011101001011100000000;
filter5[2][308] = 35'b11111011001001110011110111100000000;
filter5[2][309] = 35'b00000100010100101010100011101000000;
filter5[2][310] = 35'b11111101101011110100000101001000000;
filter5[2][311] = 35'b11111101101111110111011000100100000;
filter5[2][312] = 35'b00000100000001110111100001010000000;
filter5[2][313] = 35'b11111101110010101110110000000000000;
filter5[2][314] = 35'b11111101011000100011100110001100000;
filter5[2][315] = 35'b11111100101101001110001100010000000;
filter5[2][316] = 35'b00000011111101110010000000111100000;
filter5[2][317] = 35'b11110110000101110101000011000000000;
filter5[2][318] = 35'b00000110001010011111101010011000000;
filter5[2][319] = 35'b11110101100110110100000001000000000;
filter5[2][320] = 35'b00000000000110000011110111101111010;
filter5[2][321] = 35'b11111011100110001111111101010000000;
filter5[2][322] = 35'b11111110000010101110111010101100000;
filter5[2][323] = 35'b11111111110101110011011100010110010;
filter5[2][324] = 35'b11111100101001101010100001000100000;
filter5[2][325] = 35'b11111101000111011010110111111100000;
filter5[2][326] = 35'b11111100111111001110001100001100000;
filter5[2][327] = 35'b11111110001100111010101010111010000;
filter5[2][328] = 35'b00000001001010001001000101010000000;
filter5[2][329] = 35'b00000000110110010010000110111001000;
filter5[2][330] = 35'b00000000111111111101011011000110000;
filter5[2][331] = 35'b11111111111110010011101111101011100;
filter5[2][332] = 35'b00000000100100110011000011010101000;
filter5[2][333] = 35'b11111011000101101011111101100000000;
filter5[2][334] = 35'b11111111111111100101101000001110110;
filter5[2][335] = 35'b00000010111110101000111000110000000;
filter5[2][336] = 35'b00000001111100111110001100101100000;
filter5[2][337] = 35'b00000011000100011000100001011100000;
filter5[2][338] = 35'b00000011001111111110100011000000000;
filter5[2][339] = 35'b11111110111110100110101101000010000;
filter5[2][340] = 35'b11111111001000110010111110100000000;
filter5[2][341] = 35'b11111010111111010111011001010000000;
filter5[2][342] = 35'b00000001001110101100000000101000000;
filter5[2][343] = 35'b00000011010100101000101010011100000;
filter5[2][344] = 35'b00000100000100101101011101110000000;
filter5[2][345] = 35'b00000001111000001110101000110000000;
filter5[2][346] = 35'b00000000011010010010011010001010000;
filter5[2][347] = 35'b00000000001111011010000011100110110;
filter5[2][348] = 35'b00000010001010001100000111111000000;
filter5[2][349] = 35'b11111111110100111111110010100110110;
filter5[2][350] = 35'b00000010001011110001000000101100000;
filter5[2][351] = 35'b11111111000101111101110101011010000;
filter5[2][352] = 35'b11111111001100110011110100101100000;
filter5[2][353] = 35'b11111101111011010000101010000100000;
filter5[2][354] = 35'b11111111110110100010010000110011100;
filter5[2][355] = 35'b00000001000001010100001111000110000;
filter5[2][356] = 35'b00000000001010100110110100110011000;
filter5[2][357] = 35'b00000001010100000011111101000110000;
filter5[2][358] = 35'b00000100010111011100111011110000000;
filter5[2][359] = 35'b11111111000100010011100110110110000;
filter5[2][360] = 35'b00000011010101010101100010010000000;
filter5[2][361] = 35'b11111110100111110111011000110000000;
filter5[2][362] = 35'b11111110011110000001011111100000000;
filter5[2][363] = 35'b11111111110011011110011111111001110;
filter5[2][364] = 35'b11111011000010110011000010011000000;
filter5[2][365] = 35'b11111111110011000000101111111111100;
filter5[2][366] = 35'b00000000111100100000010110001010000;
filter5[2][367] = 35'b11111110111101100001100011010100000;
filter5[2][368] = 35'b11111111111111101110100011000000011;
filter5[2][369] = 35'b11111100000110110010111010000000000;
filter5[2][370] = 35'b11111110000000111101111011111010000;
filter5[2][371] = 35'b00000000000000001000101100100010011;
filter5[2][372] = 35'b11111101011001101111000100100000000;
filter5[2][373] = 35'b00000011101101110010111110101100000;
filter5[2][374] = 35'b11111110100100100001001001011100000;
filter5[2][375] = 35'b11111011100011111101001010100000000;
filter5[2][376] = 35'b00000001010100000001111000010100000;
filter5[2][377] = 35'b00000111110010001010010111100000000;
filter5[2][378] = 35'b00000011000101101011101010111100000;
filter5[2][379] = 35'b00000010101001001110101001100100000;
filter5[2][380] = 35'b11111011110001000111100001010000000;
filter5[2][381] = 35'b00000000011100010000110010001100100;
filter5[2][382] = 35'b00000100100011111000110111011000000;
filter5[2][383] = 35'b11111001010100011100110010001000000;
filter5[2][384] = 35'b00000010001010001100011111011100000;
filter5[2][385] = 35'b11111110100111000101011101000110000;
filter5[2][386] = 35'b11111111110001100111010101000100010;
filter5[2][387] = 35'b11111111100101001110101110011001000;
filter5[2][388] = 35'b11111101011011111000110101110100000;
filter5[2][389] = 35'b11111111000111101101001100101101000;
filter5[2][390] = 35'b00000010001010110001000110111000000;
filter5[2][391] = 35'b00000000101111000001110111100001000;
filter5[2][392] = 35'b11111110001010010010111110011010000;
filter5[2][393] = 35'b00000010001001100011011001000100000;
filter5[2][394] = 35'b00000010101011000110011110010100000;
filter5[2][395] = 35'b11111111100101101101101000011010100;
filter5[2][396] = 35'b11111101101010111101111101000000000;
filter5[2][397] = 35'b11111101010001000110100010011100000;
filter5[2][398] = 35'b11111101011010000011010010000100000;
filter5[2][399] = 35'b00000010011101011101100110100000000;
filter5[2][400] = 35'b00000001011010011000111100010100000;
filter5[2][401] = 35'b11111111000010010101000111101010000;
filter5[2][402] = 35'b00000001010000010110000001100010000;
filter5[2][403] = 35'b11111111011000011001100100101010000;
filter5[2][404] = 35'b11111101000100001101010101001100000;
filter5[2][405] = 35'b00000000110100111100010010111000000;
filter5[2][406] = 35'b11111101001001100111000101010100000;
filter5[2][407] = 35'b00000000111011111100010011001101000;
filter5[2][408] = 35'b11111110010100110111111010000010000;
filter5[2][409] = 35'b00000000111111110100001000000000000;
filter5[2][410] = 35'b00000011000010110110011100010100000;
filter5[2][411] = 35'b00000001001000010011010100101100000;
filter5[2][412] = 35'b00000001101101010111110000101010000;
filter5[2][413] = 35'b11111101101000011000010110111100000;
filter5[2][414] = 35'b11111110101011000100011111011100000;
filter5[2][415] = 35'b11111110010011100001101001001010000;
filter5[2][416] = 35'b11111110111001110110001110011100000;
filter5[2][417] = 35'b00000000000001110110101001101001011;
filter5[2][418] = 35'b11111111001110110101101010010000000;
filter5[2][419] = 35'b11111111111111001101101000001001110;
filter5[2][420] = 35'b11111110100010000110000011001000000;
filter5[2][421] = 35'b00000000100001101101100111001000000;
filter5[2][422] = 35'b00000100101001000100000100000000000;
filter5[2][423] = 35'b00000111010000000110111110001000000;
filter5[2][424] = 35'b11111110011110111111000111100100000;
filter5[2][425] = 35'b00000000110011111100001111011011000;
filter5[2][426] = 35'b00000000011110100011101100010111100;
filter5[2][427] = 35'b11111110111001001011100100101100000;
filter5[2][428] = 35'b00000000100100001110101000000100000;
filter5[2][429] = 35'b11111010100111010001010100011000000;
filter5[2][430] = 35'b00000100001011001010101011011000000;
filter5[2][431] = 35'b11111101111011001010111000011100000;
filter5[2][432] = 35'b11111111100011000101101101110101000;
filter5[2][433] = 35'b11111111010101000100110110011001000;
filter5[2][434] = 35'b11111101111000101110101101010100000;
filter5[2][435] = 35'b00000001000110100111100110110110000;
filter5[2][436] = 35'b11111111111010101011001100010001110;
filter5[2][437] = 35'b00000000101010011111111011100001000;
filter5[2][438] = 35'b00000000010101100111010101101100000;
filter5[2][439] = 35'b11111111000011100001101010110011000;
filter5[2][440] = 35'b11111110111111110010111100011010000;
filter5[2][441] = 35'b00000010100101100011001110011100000;
filter5[2][442] = 35'b00000011110001000111111001000100000;
filter5[2][443] = 35'b00000100100110001101111101001000000;
filter5[2][444] = 35'b11111101000110011111011001010100000;
filter5[2][445] = 35'b11111011011001100011100001100000000;
filter5[2][446] = 35'b00000000100110111010101110111011000;
filter5[2][447] = 35'b00000001000111101110101011000110000;
filter5[2][448] = 35'b00000011110110011100001110100100000;
filter5[2][449] = 35'b11111010100100000101001000110000000;
filter5[2][450] = 35'b00000100011101110110110010101000000;
filter5[2][451] = 35'b11111100000100101001011001110000000;
filter5[2][452] = 35'b11110101110111000001011101000000000;
filter5[2][453] = 35'b11111101110100101010110000001100000;
filter5[2][454] = 35'b00000000001110000110010000110101010;
filter5[2][455] = 35'b00000100110000011000001101100000000;
filter5[2][456] = 35'b11111010111000010100100100001000000;
filter5[2][457] = 35'b00000011111000100011010111110100000;
filter5[2][458] = 35'b00000010101010100010010001000000000;
filter5[2][459] = 35'b11110111100001001100100101000000000;
filter5[2][460] = 35'b11111001100000111111001001110000000;
filter5[2][461] = 35'b00000100111010000100001110101000000;
filter5[2][462] = 35'b00000001011110000100000110101100000;
filter5[2][463] = 35'b11111111101001110001100010010111000;
filter5[2][464] = 35'b00000000110110001111100000001101000;
filter5[2][465] = 35'b11111100010011101110001111010000000;
filter5[2][466] = 35'b11111101000101010100111000111000000;
filter5[2][467] = 35'b11111100110001011111000010101100000;
filter5[2][468] = 35'b11110011100110011001110010010000000;
filter5[2][469] = 35'b11110110110110100111001101100000000;
filter5[2][470] = 35'b00001100100100001100011101110000000;
filter5[2][471] = 35'b00000011001000001100001000001000000;
filter5[2][472] = 35'b11111111000110111001101111001100000;
filter5[2][473] = 35'b11111111010110110100110110111001000;
filter5[2][474] = 35'b11111100100111011001001000011000000;
filter5[2][475] = 35'b11111110001011100010110000000110000;
filter5[2][476] = 35'b00000011100001001101001000011100000;
filter5[2][477] = 35'b00000010011010110101111101011100000;
filter5[2][478] = 35'b00001010001011011101110101110000000;
filter5[2][479] = 35'b00000101011000010010110111000000000;
filter5[2][480] = 35'b00000011000010110110100101010000000;
filter5[2][481] = 35'b11111101110011110001111100110100000;
filter5[2][482] = 35'b11111000111000011101111000001000000;
filter5[2][483] = 35'b00000001000011001110010100111010000;
filter5[2][484] = 35'b00000001010101010111011110001000000;
filter5[2][485] = 35'b00000111010111101011001000011000000;
filter5[2][486] = 35'b00000110111000011011111111000000000;
filter5[2][487] = 35'b00000000010011110111111110010000000;
filter5[2][488] = 35'b11111101010111111010011000100100000;
filter5[2][489] = 35'b11111111101100001001110011000000000;
filter5[2][490] = 35'b11110111010111000001000001000000000;
filter5[2][491] = 35'b11111101001100100001001000101100000;
filter5[2][492] = 35'b11111111001110101100000101000110000;
filter5[2][493] = 35'b00000010001000111010110011110100000;
filter5[2][494] = 35'b00000101100100110110101110011000000;
filter5[2][495] = 35'b11111011111101110011111011001000000;
filter5[2][496] = 35'b00000010110000101001111101000100000;
filter5[2][497] = 35'b11111100101000011010000111011000000;
filter5[2][498] = 35'b11110111101110000001001000100000000;
filter5[2][499] = 35'b11111101111110101011000010001000000;
filter5[2][500] = 35'b00000000010001100010110011110111000;
filter5[2][501] = 35'b11111111110011101010010100110101000;
filter5[2][502] = 35'b11111110100001101100010000010010000;
filter5[2][503] = 35'b11111011000110001000010010010000000;
filter5[2][504] = 35'b11111110000110110110111011000010000;
filter5[2][505] = 35'b11111001101000010101111111100000000;
filter5[2][506] = 35'b11110100110111110001000111100000000;
filter5[2][507] = 35'b11111101010000011011101110100000000;
filter5[2][508] = 35'b11111101100101011001100001101100000;
filter5[2][509] = 35'b00000001001001110001110011101000000;
filter5[2][510] = 35'b00000011110000100010001110011000000;
filter5[2][511] = 35'b00000010101010101011001110100100000;
filter5[2][512] = 35'b00000001001010101101100011101000000;
filter5[2][513] = 35'b11111111000101100001100001101100000;
filter5[2][514] = 35'b11111111000100111010100000000100000;
filter5[2][515] = 35'b00000010101111110100100010111100000;
filter5[2][516] = 35'b11111011101111010001011000100000000;
filter5[2][517] = 35'b11111001110100101100110110011000000;
filter5[2][518] = 35'b11111100111000110001010000010000000;
filter5[2][519] = 35'b11111111100101100111000110101010000;
filter5[2][520] = 35'b11111111110011111111101001110001100;
filter5[2][521] = 35'b11111110110010101001100100111000000;
filter5[2][522] = 35'b00000000110011101111011001011000000;
filter5[2][523] = 35'b00000000101100111011110000100100000;
filter5[2][524] = 35'b00000011110000100101110001011100000;
filter5[2][525] = 35'b11111110110001111100000111101110000;
filter5[2][526] = 35'b11111110011100000001100001011000000;
filter5[2][527] = 35'b00000000011111101000110001010001100;
filter5[2][528] = 35'b00000001110001110011100001010110000;
filter5[2][529] = 35'b00000001001001011110000010100000000;
filter5[2][530] = 35'b00000001111001111000011011001100000;
filter5[2][531] = 35'b00000000001010111010000100001000110;
filter5[2][532] = 35'b00000000100110110010011010111010000;
filter5[2][533] = 35'b11111101111100101110100111111100000;
filter5[2][534] = 35'b11111111010001010010110110000000000;
filter5[2][535] = 35'b11111101101110001101001100010100000;
filter5[2][536] = 35'b00000001001001000000111111110000000;
filter5[2][537] = 35'b00000010110001101111001111010000000;
filter5[2][538] = 35'b00000011011001110100100000110100000;
filter5[2][539] = 35'b00000001100101110110111101011010000;
filter5[2][540] = 35'b00000001000100001001010001101010000;
filter5[2][541] = 35'b11111110000011100001001001000110000;
filter5[2][542] = 35'b11111101100110110100110100001000000;
filter5[2][543] = 35'b11111110100100110000000100101000000;
filter5[2][544] = 35'b00000000011110001001101100001011100;
filter5[2][545] = 35'b11111110010110110100000010111010000;
filter5[2][546] = 35'b11111100110011100001110011100100000;
filter5[2][547] = 35'b11111110000110000000110001010110000;
filter5[2][548] = 35'b11111111100000101110010101100100000;
filter5[2][549] = 35'b00000000110010011011111111111101000;
filter5[2][550] = 35'b00000010110110100001010010110000000;
filter5[2][551] = 35'b00000100001101110111011101011000000;
filter5[2][552] = 35'b00000010111000111011001101001100000;
filter5[2][553] = 35'b11111110001100110110111110000010000;
filter5[2][554] = 35'b11111101100111010100100000001000000;
filter5[2][555] = 35'b00000010101101001101110100111000000;
filter5[2][556] = 35'b00000010110011000001110001111000000;
filter5[2][557] = 35'b00000010101000011101100111101000000;
filter5[2][558] = 35'b00000000111101000011101111010000000;
filter5[2][559] = 35'b11111101011101110011111001011000000;
filter5[2][560] = 35'b00000000011001000010000001111110000;
filter5[2][561] = 35'b00000000010001001000101011011011100;
filter5[2][562] = 35'b11111110110001111010101001111100000;
filter5[2][563] = 35'b11111111100110101111100110111011000;
filter5[2][564] = 35'b11111110110010000010111101100010000;
filter5[2][565] = 35'b11111101010110111110010001001000000;
filter5[2][566] = 35'b11111101110010111110010010101000000;
filter5[2][567] = 35'b11111101101100101011000011001100000;
filter5[2][568] = 35'b00000001101110011001011000100110000;
filter5[2][569] = 35'b00000000100011100011010001100101000;
filter5[2][570] = 35'b00000010100000001010101001000100000;
filter5[2][571] = 35'b00000001011011000001011001001010000;
filter5[2][572] = 35'b11111111110111011001011001000111010;
filter5[2][573] = 35'b00000000100001000010100011100000000;
filter5[2][574] = 35'b11111111011001101011101011100111000;
filter5[2][575] = 35'b11111111001010010010110000100011000;
filter5[2][576] = 35'b00000001101101110010101100110000000;
filter5[2][577] = 35'b11111111111011001011101010100111010;
filter5[2][578] = 35'b00000011110000101110011001101000000;
filter5[2][579] = 35'b00000101000111011001100111000000000;
filter5[2][580] = 35'b11111111110000111000101100110001110;
filter5[2][581] = 35'b11111110001010010110111000011000000;
filter5[2][582] = 35'b11111111010111110111000100010111000;
filter5[2][583] = 35'b00000000110010000010010011010110000;
filter5[2][584] = 35'b00000000100010110101111001110100000;
filter5[2][585] = 35'b00000000110111000000100110101010000;
filter5[2][586] = 35'b00000001111011110101101010110010000;
filter5[2][587] = 35'b11111111101000001111111010100011000;
filter5[2][588] = 35'b11111111111100011111111110111010101;
filter5[2][589] = 35'b11111011010010011000111001011000000;
filter5[2][590] = 35'b11111110001110110110101010101100000;
filter5[2][591] = 35'b00000000010001011101100110111100000;
filter5[2][592] = 35'b00000010110010001010011001000000000;
filter5[2][593] = 35'b11111101101100110110010011100100000;
filter5[2][594] = 35'b00000000111110111001001010101101000;
filter5[2][595] = 35'b11111100010101110110100010011000000;
filter5[2][596] = 35'b00000001101010111111111100100100000;
filter5[2][597] = 35'b11111110011100110110010110110110000;
filter5[2][598] = 35'b11111101011110100111110101100000000;
filter5[2][599] = 35'b11111100101001110111111000110100000;
filter5[2][600] = 35'b00000000100111001001100100000100000;
filter5[2][601] = 35'b00000010010100111010101001111100000;
filter5[2][602] = 35'b11111100111110001000000011100100000;
filter5[2][603] = 35'b00000001000100000100101001101100000;
filter5[2][604] = 35'b00000111100101010101001101100000000;
filter5[2][605] = 35'b00000000100011101101101100010110000;
filter5[2][606] = 35'b00000000111011000010101100101101000;
filter5[2][607] = 35'b11111111111010010101000111010000110;
filter5[2][608] = 35'b00000100000110100110000110101000000;
filter5[2][609] = 35'b00000011011010111100110101001000000;
filter5[2][610] = 35'b11111111111001101011100100000011001;
filter5[2][611] = 35'b11111101111001101000101100001000000;
filter5[2][612] = 35'b00000010000010011001011001111000000;
filter5[2][613] = 35'b11111111000111101000010001110111000;
filter5[2][614] = 35'b00000011001111001001100000010100000;
filter5[2][615] = 35'b00000001111111000110011010010100000;
filter5[2][616] = 35'b00000000011010101101001010110110000;
filter5[2][617] = 35'b00000011000011110101101111011000000;
filter5[2][618] = 35'b11111011011000000101011111001000000;
filter5[2][619] = 35'b11111011011001100000011011001000000;
filter5[2][620] = 35'b11111011111100010101111100100000000;
filter5[2][621] = 35'b00000000001111111101000011010000100;
filter5[2][622] = 35'b00000000110111111001101110110111000;
filter5[2][623] = 35'b11111101011111001001011011111000000;
filter5[2][624] = 35'b11111111110001001110011010010011000;
filter5[2][625] = 35'b00000101000100001110111111101000000;
filter5[2][626] = 35'b11111101101111110010110001011000000;
filter5[2][627] = 35'b00000010010111000100000000010000000;
filter5[2][628] = 35'b00000000100010101000001100011011000;
filter5[2][629] = 35'b11111010100010010011110000001000000;
filter5[2][630] = 35'b11111110000110101111000111101110000;
filter5[2][631] = 35'b11111110110100101000010010011010000;
filter5[2][632] = 35'b00000001011011100110011011000100000;
filter5[2][633] = 35'b00000011001010000110100110000000000;
filter5[2][634] = 35'b00000100011000000010011100001000000;
filter5[2][635] = 35'b00000001001101101110010001010100000;
filter5[2][636] = 35'b00000000001010101010101101000011110;
filter5[2][637] = 35'b00000010000110011110010011110100000;
filter5[2][638] = 35'b11111110011011100100101111100110000;
filter5[2][639] = 35'b00000001100010101011111100010100000;
filter5[2][640] = 35'b11111110110101010100111110001010000;
filter5[2][641] = 35'b11110011111100111001101011100000000;
filter5[2][642] = 35'b11111111000010010000010011100010000;
filter5[2][643] = 35'b11111100000001110010110011101000000;
filter5[2][644] = 35'b11111001110101100111100100000000000;
filter5[2][645] = 35'b11111111010000100011000111010101000;
filter5[2][646] = 35'b00000001101101001001110001010000000;
filter5[2][647] = 35'b11111101111001101011111100110000000;
filter5[2][648] = 35'b00000011101101101100000001110000000;
filter5[2][649] = 35'b00000001010010000001110001101110000;
filter5[2][650] = 35'b00000010111101111011101010010000000;
filter5[2][651] = 35'b11111001110000011111100100110000000;
filter5[2][652] = 35'b11111010000011011100111010111000000;
filter5[2][653] = 35'b11111110101110100001100010001010000;
filter5[2][654] = 35'b00000000000001001001001101010011100;
filter5[2][655] = 35'b00000011000100110110000011001100000;
filter5[2][656] = 35'b00000000001100111001011101000001000;
filter5[2][657] = 35'b11111110001001010101010000000110000;
filter5[2][658] = 35'b00000011000010100110010111001000000;
filter5[2][659] = 35'b11111011011000101110011111100000000;
filter5[2][660] = 35'b00000011110011100100010100011000000;
filter5[2][661] = 35'b11111000101100110110110101111000000;
filter5[2][662] = 35'b11111101111010110001100101111100000;
filter5[2][663] = 35'b11111010101000010110001111110000000;
filter5[2][664] = 35'b00000000001011110111110110011011100;
filter5[2][665] = 35'b00000011011000110111100100011000000;
filter5[2][666] = 35'b00000001111100100010110110011010000;
filter5[2][667] = 35'b11111111110001101000101011000101010;
filter5[2][668] = 35'b11111011101110101110110101011000000;
filter5[2][669] = 35'b11111010110110000000001100000000000;
filter5[2][670] = 35'b11111110110100011100001110010100000;
filter5[2][671] = 35'b00000001000010111100010010001110000;
filter5[2][672] = 35'b00000010101100111010110011000100000;
filter5[2][673] = 35'b00000010011010100001011100011000000;
filter5[2][674] = 35'b11111111001001000101011111011000000;
filter5[2][675] = 35'b00000001010001110000001110000010000;
filter5[2][676] = 35'b00000101100000010010001110101000000;
filter5[2][677] = 35'b00000001101101011011011001101100000;
filter5[2][678] = 35'b00001000011100000111001110100000000;
filter5[2][679] = 35'b00000010000001010100010011110100000;
filter5[2][680] = 35'b11111111110001000000010111011000000;
filter5[2][681] = 35'b00000010110001100011011000100100000;
filter5[2][682] = 35'b11111011111010101110100011111000000;
filter5[2][683] = 35'b00000001111100111110111000011100000;
filter5[2][684] = 35'b00000010001001010110100000111000000;
filter5[2][685] = 35'b00000011011011111011011000100100000;
filter5[2][686] = 35'b00000011000010111110101000010100000;
filter5[2][687] = 35'b11111100000111100100000000001100000;
filter5[2][688] = 35'b00000011101010101100111011011100000;
filter5[2][689] = 35'b00000001010110011111011011000100000;
filter5[2][690] = 35'b00000000100000000010110110001110000;
filter5[2][691] = 35'b11111011000110100101011111000000000;
filter5[2][692] = 35'b11111110000010100100010010100000000;
filter5[2][693] = 35'b11111110010011111001010011001010000;
filter5[2][694] = 35'b11111111101100100011001100000100000;
filter5[2][695] = 35'b11111011001111111101110001000000000;
filter5[2][696] = 35'b11111011011110110001100011110000000;
filter5[2][697] = 35'b11111101110011010111011000101100000;
filter5[2][698] = 35'b00000001111000011111001111111010000;
filter5[2][699] = 35'b00000000110001110101110111001110000;
filter5[2][700] = 35'b11111010111110011000000011011000000;
filter5[2][701] = 35'b11111111101010100011001011100111000;
filter5[2][702] = 35'b00000010110000111010001001100000000;
filter5[2][703] = 35'b00000010110011000110000000001000000;
filter5[2][704] = 35'b11111110100101111011101110001000000;
filter5[2][705] = 35'b00000000001001110111100000011000010;
filter5[2][706] = 35'b11111111000100010101000001010001000;
filter5[2][707] = 35'b11111110001111100010011100101100000;
filter5[2][708] = 35'b00000000101001100100010101001101000;
filter5[2][709] = 35'b11111101011110000111111111100000000;
filter5[2][710] = 35'b11111111100010010011010010100110100;
filter5[2][711] = 35'b00000000000110110011111011010010010;
filter5[2][712] = 35'b11111111010001110111001011011101000;
filter5[2][713] = 35'b11111101011111011010110100111000000;
filter5[2][714] = 35'b00000000011111000110100111011010000;
filter5[2][715] = 35'b11111111010000001011000011010100000;
filter5[2][716] = 35'b00000001011110110001011101001110000;
filter5[2][717] = 35'b11111101011101000101111011000100000;
filter5[2][718] = 35'b11111110111111000101111010000110000;
filter5[2][719] = 35'b00000010110101111000000110111000000;
filter5[2][720] = 35'b00000000011100101101110011011100000;
filter5[2][721] = 35'b00000000110011000000110001100010000;
filter5[2][722] = 35'b11111010100110001100000111000000000;
filter5[2][723] = 35'b00000001100101001101100110010000000;
filter5[2][724] = 35'b00000000000000100000011100010000110;
filter5[2][725] = 35'b11111100111001110111111000100100000;
filter5[2][726] = 35'b00000000000001011111101100011000001;
filter5[2][727] = 35'b00000100000001111100101000000000000;
filter5[2][728] = 35'b11111111011101111011010000110111000;
filter5[2][729] = 35'b11111111110001010000110100011111110;
filter5[2][730] = 35'b11111110011000110110000010010010000;
filter5[2][731] = 35'b00000000000101111101111100000101101;
filter5[2][732] = 35'b11111011010111101010100000100000000;
filter5[2][733] = 35'b00000010101111000100010111111100000;
filter5[2][734] = 35'b00000100100100011111111000100000000;
filter5[2][735] = 35'b00000010001001110011001100001000000;
filter5[2][736] = 35'b00000000001101101000111011011100010;
filter5[2][737] = 35'b11111111110010010111100010000010010;
filter5[2][738] = 35'b11111011001011100000001100100000000;
filter5[2][739] = 35'b00000000001101001110110000001111100;
filter5[2][740] = 35'b00000001010110000001110011000000000;
filter5[2][741] = 35'b00000101110011011011101010011000000;
filter5[2][742] = 35'b00000011011001111100111011111000000;
filter5[2][743] = 35'b11111100110110001110000101101100000;
filter5[2][744] = 35'b11111110010101000110001010000010000;
filter5[2][745] = 35'b11111100011110100000001110001000000;
filter5[2][746] = 35'b00000000100110010111000110011011000;
filter5[2][747] = 35'b11111010111011011101101101000000000;
filter5[2][748] = 35'b11111100111010110011110111111100000;
filter5[2][749] = 35'b00000001110000101001111110100010000;
filter5[2][750] = 35'b00000100001011110000111110111000000;
filter5[2][751] = 35'b11111011111010100100100111110000000;
filter5[2][752] = 35'b11111110000000100111111001110110000;
filter5[2][753] = 35'b00000000100011100010001001001101000;
filter5[2][754] = 35'b11111101000100100000010110001000000;
filter5[2][755] = 35'b11111110111100010110001010110110000;
filter5[2][756] = 35'b11111101100000110011100010000000000;
filter5[2][757] = 35'b11111111000111110101100001101001000;
filter5[2][758] = 35'b11111010111111000011011100010000000;
filter5[2][759] = 35'b11111011000110011101001000100000000;
filter5[2][760] = 35'b11111101011110101000100000001000000;
filter5[2][761] = 35'b11111111100001111101111111010011000;
filter5[2][762] = 35'b00000001110000001000110101010100000;
filter5[2][763] = 35'b00000010000011011000111010110100000;
filter5[2][764] = 35'b11111110001110000101000001101010000;
filter5[2][765] = 35'b11111100000100011101101001111100000;
filter5[2][766] = 35'b00000000111000110100111011111110000;
filter5[2][767] = 35'b11111100110001011101001010101000000;
filter5[2][768] = 35'b11111011100110111101100110000000000;
filter5[2][769] = 35'b00000000101010101001100000011100000;
filter5[2][770] = 35'b11111110110000001001101001011000000;
filter5[2][771] = 35'b11111101011000110010110111011100000;
filter5[2][772] = 35'b11111100100010111010011010100000000;
filter5[2][773] = 35'b00000000110000100010010010010111000;
filter5[2][774] = 35'b00000001011000110110000000100100000;
filter5[2][775] = 35'b00000010001110111111101001101100000;
filter5[2][776] = 35'b11111110010011000001110000101100000;
filter5[2][777] = 35'b00000000010011010110111110100001000;
filter5[2][778] = 35'b11111100010001000111000101010000000;
filter5[2][779] = 35'b00000000100010001111000111101110000;
filter5[2][780] = 35'b11111100110001100011111001111100000;
filter5[2][781] = 35'b11111001001010110100100110000000000;
filter5[2][782] = 35'b00000101011110000000101000001000000;
filter5[2][783] = 35'b11111111001111001100000011001010000;
filter5[2][784] = 35'b00000000101101110000001100010111000;
filter5[2][785] = 35'b00000000010100111100001011110111100;
filter5[2][786] = 35'b11111110110001001110011001011010000;
filter5[2][787] = 35'b11111110000001110111100001010100000;
filter5[2][788] = 35'b11111100011011001110111100011100000;
filter5[2][789] = 35'b00000011010000101000010000000000000;
filter5[2][790] = 35'b00001000001001001000101010010000000;
filter5[2][791] = 35'b00000010111110011001000100000100000;
filter5[2][792] = 35'b00000000000001100000101001010101100;
filter5[2][793] = 35'b00000000001001010010001110010000010;
filter5[2][794] = 35'b11111100101100001110010111011100000;
filter5[2][795] = 35'b00000010110010110110001000000000000;
filter5[2][796] = 35'b11111111101001010011110101000111000;
filter5[2][797] = 35'b00000110010010100011100111111000000;
filter5[2][798] = 35'b00000101000010000100000111010000000;
filter5[2][799] = 35'b00000011100110111010001100100100000;
filter5[2][800] = 35'b11111110001111111001101001110010000;
filter5[2][801] = 35'b11111100100110011110110000100100000;
filter5[2][802] = 35'b11111100110101110110011110000000000;
filter5[2][803] = 35'b00000000011101110000110101000010100;
filter5[2][804] = 35'b11111110100111000011001111010000000;
filter5[2][805] = 35'b00001010100101001110110101000000000;
filter5[2][806] = 35'b00000110111111000101001100110000000;
filter5[2][807] = 35'b00000111011110001011111001101000000;
filter5[2][808] = 35'b11111101011010111001100010101100000;
filter5[2][809] = 35'b11111110100000010011110101110110000;
filter5[2][810] = 35'b11111101101111111111011101111000000;
filter5[2][811] = 35'b11111111101000111101000011100001100;
filter5[2][812] = 35'b00000001100101001101001000101110000;
filter5[2][813] = 35'b00000101100011000010101110010000000;
filter5[2][814] = 35'b00000101010011111011111001100000000;
filter5[2][815] = 35'b11111111011110111110011000001000000;
filter5[2][816] = 35'b00000001010000010101100101111010000;
filter5[2][817] = 35'b11111111100011001110001100110110100;
filter5[2][818] = 35'b11111110010001110111011000010110000;
filter5[2][819] = 35'b11110110101100001101000011110000000;
filter5[2][820] = 35'b11111101010011001100101001011100000;
filter5[2][821] = 35'b11111111010101100110000010100010000;
filter5[2][822] = 35'b11111110001000010011100100101000000;
filter5[2][823] = 35'b11111101011100001001101111110100000;
filter5[2][824] = 35'b00000100000100000100010001010000000;
filter5[2][825] = 35'b00000101111101011111110100111000000;
filter5[2][826] = 35'b11111101111010100101001000101100000;
filter5[2][827] = 35'b00000000111100110011111111011000000;
filter5[2][828] = 35'b11111010000100000000110101001000000;
filter5[2][829] = 35'b11111111011101000000010110110010000;
filter5[2][830] = 35'b00000000110010010000010110101001000;
filter5[2][831] = 35'b11111101101010111101011000000100000;
filter5[2][832] = 35'b00000000101011110000011010001011000;
filter5[2][833] = 35'b00000000000000000000100011001101011;
filter5[2][834] = 35'b11111111111110010001111011000110000;
filter5[2][835] = 35'b00000000001111011011110101011011100;
filter5[2][836] = 35'b11111110110101100011111111011110000;
filter5[2][837] = 35'b11111111011001001000101101010100000;
filter5[2][838] = 35'b11111110111100110110100010000000000;
filter5[2][839] = 35'b11111111010000110001001101101011000;
filter5[2][840] = 35'b11111111010000001010110101001001000;
filter5[2][841] = 35'b11111111001101010010101001000001000;
filter5[2][842] = 35'b00000001001010011010101001100000000;
filter5[2][843] = 35'b11111111001100010010101110001111000;
filter5[2][844] = 35'b11111101101011001111100011000100000;
filter5[2][845] = 35'b00000010000110110010110110100100000;
filter5[2][846] = 35'b11111111100101100100001100011110000;
filter5[2][847] = 35'b11111110001101110110101110010010000;
filter5[2][848] = 35'b00000000101110000011110011100010000;
filter5[2][849] = 35'b00000001001000000101101010010000000;
filter5[2][850] = 35'b00000000101101100111001111101111000;
filter5[2][851] = 35'b00000100010011010001100100100000000;
filter5[2][852] = 35'b11111111100111011010100101001111000;
filter5[2][853] = 35'b11111000100001010000011010100000000;
filter5[2][854] = 35'b00000000100101011011100111111000000;
filter5[2][855] = 35'b00000101111101101100011010111000000;
filter5[2][856] = 35'b00000001010000000110111011100100000;
filter5[2][857] = 35'b11111100110101110100011001110000000;
filter5[2][858] = 35'b11110110110001001100111011010000000;
filter5[2][859] = 35'b00000110001100110110110011010000000;
filter5[2][860] = 35'b11111011111100100101100011100000000;
filter5[2][861] = 35'b00000100101001000010001111001000000;
filter5[2][862] = 35'b00000000101100000001101110101001000;
filter5[2][863] = 35'b00000100001000111100001111110000000;
filter5[2][864] = 35'b11111110001010000000000010011100000;
filter5[2][865] = 35'b11111010101110111010100001000000000;
filter5[2][866] = 35'b11111110100101001100010100000100000;
filter5[2][867] = 35'b00000001000110100100111111011110000;
filter5[2][868] = 35'b11111100010001011101001100110100000;
filter5[2][869] = 35'b00000010010001000111101111001000000;
filter5[2][870] = 35'b11111111100010010010010111100111000;
filter5[2][871] = 35'b11111001100010001000111111001000000;
filter5[2][872] = 35'b00000001101101000000110010000000000;
filter5[2][873] = 35'b11111010101110011001010000110000000;
filter5[2][874] = 35'b11111111110111000000101001011001010;
filter5[2][875] = 35'b11111101011101000001000100100100000;
filter5[2][876] = 35'b00000001110010101111101111001100000;
filter5[2][877] = 35'b00000100000110010011001011010000000;
filter5[2][878] = 35'b11111101110001000001110001011000000;
filter5[2][879] = 35'b00000100001000001011000110010000000;
filter5[2][880] = 35'b11111111111101101111100101101011100;
filter5[2][881] = 35'b11111101000100001110110010001100000;
filter5[2][882] = 35'b11111100011000010011000100101100000;
filter5[2][883] = 35'b11111001011101111110110100011000000;
filter5[2][884] = 35'b00000000110100011000011111000111000;
filter5[2][885] = 35'b11111111101010001000100000001000100;
filter5[2][886] = 35'b11111110000111111010111000000000000;
filter5[2][887] = 35'b11111101001011010001111001111100000;
filter5[2][888] = 35'b11111101100111011010101001010000000;
filter5[2][889] = 35'b11111100111110010101101010111000000;
filter5[2][890] = 35'b11111101011010010101111101100000000;
filter5[2][891] = 35'b11111110010110101111011100000010000;
filter5[2][892] = 35'b11111101001100000000110111010100000;
filter5[2][893] = 35'b00000011011000001100100111011000000;
filter5[2][894] = 35'b11111000010111100111000100001000000;
filter5[2][895] = 35'b11111110110000000001111110100110000;
filter5[2][896] = 35'b11111101001000000010111010100000000;
filter5[2][897] = 35'b11111010011010011000111001010000000;
filter5[2][898] = 35'b00000010000000011100001100000100000;
filter5[2][899] = 35'b00000000110100001110001101101110000;
filter5[2][900] = 35'b11111110111100011011101100111010000;
filter5[2][901] = 35'b11111101001110011110110010001000000;
filter5[2][902] = 35'b11111001111110111000110010000000000;
filter5[2][903] = 35'b00000010101010010011010100100000000;
filter5[2][904] = 35'b11111101100111011110110101110000000;
filter5[2][905] = 35'b11110110110110101111000001010000000;
filter5[2][906] = 35'b11111010101110110001000001110000000;
filter5[2][907] = 35'b00000000000101100010111000111000011;
filter5[2][908] = 35'b00000010011010111111110011000100000;
filter5[2][909] = 35'b11111010010101111111111100101000000;
filter5[2][910] = 35'b11111001010010010110100110101000000;
filter5[2][911] = 35'b11111011100101110011101110001000000;
filter5[2][912] = 35'b00000001011001101010001100111010000;
filter5[2][913] = 35'b11111000011011011010101111010000000;
filter5[2][914] = 35'b11110111110111111011101001000000000;
filter5[2][915] = 35'b00000000110100100111101000111000000;
filter5[2][916] = 35'b00000001001100101010001011001110000;
filter5[2][917] = 35'b11111110011001100110110010111010000;
filter5[2][918] = 35'b00000010111011011001011001011100000;
filter5[2][919] = 35'b00001100001110010000010001010000000;
filter5[2][920] = 35'b00000010110100010001000100100100000;
filter5[2][921] = 35'b11101111100100001000110100000000000;
filter5[2][922] = 35'b11111000110000111111001011001000000;
filter5[2][923] = 35'b00000000110110101100011100010111000;
filter5[2][924] = 35'b11111100101111110010001001101000000;
filter5[2][925] = 35'b00000010011110000111110010011100000;
filter5[2][926] = 35'b00000011000100100001010100101100000;
filter5[2][927] = 35'b00000000101100011111100111111011000;
filter5[2][928] = 35'b11111101000101011000010001000100000;
filter5[2][929] = 35'b11110110100110110100000001110000000;
filter5[2][930] = 35'b11111100111000100010000110100000000;
filter5[2][931] = 35'b00000001000010001000100100110100000;
filter5[2][932] = 35'b00000000101001101000111100000110000;
filter5[2][933] = 35'b00000100000001011001011011110000000;
filter5[2][934] = 35'b00000010010011001000001011100000000;
filter5[2][935] = 35'b11110100110001000001101110000000000;
filter5[2][936] = 35'b00000011101101101110010011110000000;
filter5[2][937] = 35'b11110011100000100110011011100000000;
filter5[2][938] = 35'b00000001010101010100110010110100000;
filter5[2][939] = 35'b11111010100001000000111101010000000;
filter5[2][940] = 35'b11111011010100011011000001000000000;
filter5[2][941] = 35'b00000001011001100010000010011010000;
filter5[2][942] = 35'b11111001110101010000000001111000000;
filter5[2][943] = 35'b11110110001010100110100011010000000;
filter5[2][944] = 35'b11111011010001100001011001110000000;
filter5[2][945] = 35'b11111110010100100001000111100110000;
filter5[2][946] = 35'b11111110100001111011111111110000000;
filter5[2][947] = 35'b11111100110110011000011100101100000;
filter5[2][948] = 35'b11110111101110011011110111100000000;
filter5[2][949] = 35'b00000101010110110001111010101000000;
filter5[2][950] = 35'b00000010111011100011101010111000000;
filter5[2][951] = 35'b11110101110010101101001001100000000;
filter5[2][952] = 35'b11111110001000100011101001011000000;
filter5[2][953] = 35'b00000101010000000010111010100000000;
filter5[2][954] = 35'b00000010000100101100000000110100000;
filter5[2][955] = 35'b11111010110011111011100101111000000;
filter5[2][956] = 35'b00000010110010011110101000111100000;
filter5[2][957] = 35'b11110010011110110100010011100000000;
filter5[2][958] = 35'b11100111100110111100010111100000000;
filter5[2][959] = 35'b11110110011000000010011101100000000;
filter5[2][960] = 35'b00000010011101011010101010100100000;
filter5[2][961] = 35'b11111110011100110010011010101100000;
filter5[2][962] = 35'b00000011010110001111011111001100000;
filter5[2][963] = 35'b11111111001110101111110110101100000;
filter5[2][964] = 35'b11111001000000100110000000111000000;
filter5[2][965] = 35'b11111100000001011101001111111100000;
filter5[2][966] = 35'b11111011100000010010111110011000000;
filter5[2][967] = 35'b11111111110110110000011000011100110;
filter5[2][968] = 35'b11111110011101110111000010101110000;
filter5[2][969] = 35'b00000010011111110000010110011100000;
filter5[2][970] = 35'b11111110010001100100010100010010000;
filter5[2][971] = 35'b11111101110010101110100101000000000;
filter5[2][972] = 35'b00000010111011101010110010100100000;
filter5[2][973] = 35'b11111110100011001001110111000000000;
filter5[2][974] = 35'b00000000000110001110101011100110000;
filter5[2][975] = 35'b00000000110011001011110110100101000;
filter5[2][976] = 35'b00000010000011100000010101000100000;
filter5[2][977] = 35'b11111111000101001101010001000011000;
filter5[2][978] = 35'b11111010010011000001000011001000000;
filter5[2][979] = 35'b00000000111000101101011010111000000;
filter5[2][980] = 35'b00000000110110100001101011011101000;
filter5[2][981] = 35'b11111111000110000101100100000100000;
filter5[2][982] = 35'b00000001001100110100010010000110000;
filter5[2][983] = 35'b00000011001011101110011011000100000;
filter5[2][984] = 35'b11111100101111011110001101011000000;
filter5[2][985] = 35'b11111000100110010001101000101000000;
filter5[2][986] = 35'b11111101011010011111011001111100000;
filter5[2][987] = 35'b11111100100110101011101000110000000;
filter5[2][988] = 35'b00000000010100110100111110001111100;
filter5[2][989] = 35'b00000010011101000111010000100100000;
filter5[2][990] = 35'b00000000000100011100000100011010010;
filter5[2][991] = 35'b11111101110011011010011111111000000;
filter5[2][992] = 35'b11111111010010000001001111100011000;
filter5[2][993] = 35'b11111010111010000101000111110000000;
filter5[2][994] = 35'b11110101011100001011011010110000000;
filter5[2][995] = 35'b11110111100010100010010100110000000;
filter5[2][996] = 35'b00000101100100011101000011101000000;
filter5[2][997] = 35'b00000001111001111011000110101010000;
filter5[2][998] = 35'b11111100111111010110111100100100000;
filter5[2][999] = 35'b00000001110111010010001110101010000;
filter5[2][1000] = 35'b00000001101000110110010011000110000;
filter5[2][1001] = 35'b00000010001011101110111111111100000;
filter5[2][1002] = 35'b11111000111111111000110000100000000;
filter5[2][1003] = 35'b11110101101000010110101011000000000;
filter5[2][1004] = 35'b11111011110010100100110110111000000;
filter5[2][1005] = 35'b11111011101110110011010001011000000;
filter5[2][1006] = 35'b11111011001110101101110011010000000;
filter5[2][1007] = 35'b00000111100101011000111101111000000;
filter5[2][1008] = 35'b11111101101111101011110111011100000;
filter5[2][1009] = 35'b11111110001111111011000101101110000;
filter5[2][1010] = 35'b11111001000011011111111101101000000;
filter5[2][1011] = 35'b11110010110100010100011011100000000;
filter5[2][1012] = 35'b11101101010011111110101100100000000;
filter5[2][1013] = 35'b11101000111011100010010111100000000;
filter5[2][1014] = 35'b11110100011100101101001110000000000;
filter5[2][1015] = 35'b11111110101100100111000011011100000;
filter5[2][1016] = 35'b11111111100110111101110001101011000;
filter5[2][1017] = 35'b11111101000100111100101011100000000;
filter5[2][1018] = 35'b00000101010010011010010010010000000;
filter5[2][1019] = 35'b11111111000100101011111100110010000;
filter5[2][1020] = 35'b00000000110011001100111001111010000;
filter5[2][1021] = 35'b11111111000101001100010011011000000;
filter5[2][1022] = 35'b11111100011110110001100010011000000;
filter5[2][1023] = 35'b00000010011001101100110100100100000;
filter5[3][0] = 35'b11111001100001001000000110101000000;
filter5[3][1] = 35'b11110110010011001001111000000000000;
filter5[3][2] = 35'b11111111011111101111101001110011000;
filter5[3][3] = 35'b00000010100000111010110110001000000;
filter5[3][4] = 35'b00000011110110101110010100000000000;
filter5[3][5] = 35'b11111000110100011010010101111000000;
filter5[3][6] = 35'b11111011111100011110100000010000000;
filter5[3][7] = 35'b11110000010001101001011000010000000;
filter5[3][8] = 35'b11111110100111001110001010111000000;
filter5[3][9] = 35'b00000101100011001010010101011000000;
filter5[3][10] = 35'b00000101011011001010101101111000000;
filter5[3][11] = 35'b00000011100110001110001011100100000;
filter5[3][12] = 35'b00000010001001100110101110101000000;
filter5[3][13] = 35'b00000000010101101110011010101110100;
filter5[3][14] = 35'b11111111000111010101111101101001000;
filter5[3][15] = 35'b11111110101111100001110001101010000;
filter5[3][16] = 35'b00000000110110110111101011001001000;
filter5[3][17] = 35'b00000011011101111011101010110100000;
filter5[3][18] = 35'b00000000100000111000011001110111000;
filter5[3][19] = 35'b11111011100011011111001100001000000;
filter5[3][20] = 35'b11111111101101100111111010101001000;
filter5[3][21] = 35'b11111110101100011001101100001100000;
filter5[3][22] = 35'b00000111010111110010000101011000000;
filter5[3][23] = 35'b00000000000101111111100111111001101;
filter5[3][24] = 35'b11111110101100000011001110011000000;
filter5[3][25] = 35'b00000011011101011000010100010000000;
filter5[3][26] = 35'b00000101101000111100111011010000000;
filter5[3][27] = 35'b11111110001010011101101110110100000;
filter5[3][28] = 35'b11111101001011011100100010001100000;
filter5[3][29] = 35'b11110111011100101100000001100000000;
filter5[3][30] = 35'b00000001011111011100001111110010000;
filter5[3][31] = 35'b00000001111001010111011111111110000;
filter5[3][32] = 35'b00000010011111010110110110000000000;
filter5[3][33] = 35'b00000011010101100010010111010100000;
filter5[3][34] = 35'b11111010010000111001100101000000000;
filter5[3][35] = 35'b11111011101011110111100010111000000;
filter5[3][36] = 35'b11111010100111110010100100011000000;
filter5[3][37] = 35'b00000010011101000101001011011000000;
filter5[3][38] = 35'b00000011111011000111000100001000000;
filter5[3][39] = 35'b00000010001100111101110011011100000;
filter5[3][40] = 35'b00000100010101100001001101101000000;
filter5[3][41] = 35'b00000010110100001101111010100100000;
filter5[3][42] = 35'b11111010011101010110010101111000000;
filter5[3][43] = 35'b11111011110010000000011010100000000;
filter5[3][44] = 35'b11111110001110011111000011111110000;
filter5[3][45] = 35'b11111100010001100000110001100100000;
filter5[3][46] = 35'b00000011100001000111101100110100000;
filter5[3][47] = 35'b11111111010010111101110110110110000;
filter5[3][48] = 35'b00000000000110001111100000101011100;
filter5[3][49] = 35'b11111110111000010001101010100010000;
filter5[3][50] = 35'b00000001111101001101100011011010000;
filter5[3][51] = 35'b11111101100100101110111000010100000;
filter5[3][52] = 35'b11111110000111101111011101110000000;
filter5[3][53] = 35'b00000000111110010110101110001000000;
filter5[3][54] = 35'b00000101111000110000010110010000000;
filter5[3][55] = 35'b11111110000001000000001000010110000;
filter5[3][56] = 35'b11111101110111101100000101111000000;
filter5[3][57] = 35'b00000100001011000100100111111000000;
filter5[3][58] = 35'b00000000110100000110110110011111000;
filter5[3][59] = 35'b00000000000011000000101001010001110;
filter5[3][60] = 35'b00000001111011000001100100000010000;
filter5[3][61] = 35'b00000010110100010110111101101000000;
filter5[3][62] = 35'b00000010111011100001010101000100000;
filter5[3][63] = 35'b11111110011111101100000101111100000;
filter5[3][64] = 35'b11111101101110100010111011110000000;
filter5[3][65] = 35'b11111011000010010011001010111000000;
filter5[3][66] = 35'b11111111010111110001001010000010000;
filter5[3][67] = 35'b00000011100110110010111100011100000;
filter5[3][68] = 35'b00000010110101000101110001011000000;
filter5[3][69] = 35'b00000010011111011000000110000100000;
filter5[3][70] = 35'b11111100100110000001001101101000000;
filter5[3][71] = 35'b11110100110111010110111101100000000;
filter5[3][72] = 35'b11111101110001110001100111101100000;
filter5[3][73] = 35'b00000100100010110101110111001000000;
filter5[3][74] = 35'b00000010110100100000111011010000000;
filter5[3][75] = 35'b00000000101110000110101110000001000;
filter5[3][76] = 35'b00000001101101000100011011100100000;
filter5[3][77] = 35'b00000010011110100001110001111000000;
filter5[3][78] = 35'b11111101100110011111110111001000000;
filter5[3][79] = 35'b00000110101011100100000111001000000;
filter5[3][80] = 35'b00000100011100000000010100000000000;
filter5[3][81] = 35'b00000010011110011011101110011100000;
filter5[3][82] = 35'b00000001100100110010110111011000000;
filter5[3][83] = 35'b11111100100011000110110011010000000;
filter5[3][84] = 35'b11111110110011010111100100010100000;
filter5[3][85] = 35'b00000001001001101000111000110110000;
filter5[3][86] = 35'b11111111101001010100001111100110000;
filter5[3][87] = 35'b11111101100000101100000101000000000;
filter5[3][88] = 35'b11111101101011101101010100000000000;
filter5[3][89] = 35'b00000010111100001000011110011100000;
filter5[3][90] = 35'b00000011100000001010000000000100000;
filter5[3][91] = 35'b11111111111011110110011011000010001;
filter5[3][92] = 35'b00000000000101010010110101011001000;
filter5[3][93] = 35'b00000000101110010101001101001000000;
filter5[3][94] = 35'b11111111101111010000000010110110000;
filter5[3][95] = 35'b11111110110110101011001111001000000;
filter5[3][96] = 35'b00000011010001011110011110001100000;
filter5[3][97] = 35'b00000001011001100010011011001010000;
filter5[3][98] = 35'b11111011100011011110110011010000000;
filter5[3][99] = 35'b11111111001001110001101001110000000;
filter5[3][100] = 35'b11111111010001111001010001110010000;
filter5[3][101] = 35'b00000000000010100111100000001010100;
filter5[3][102] = 35'b11111011010100000000000111010000000;
filter5[3][103] = 35'b11111111111001100000010111010010001;
filter5[3][104] = 35'b00000101111001000010010011111000000;
filter5[3][105] = 35'b00000001000010000100101000010110000;
filter5[3][106] = 35'b11111110010101010000011110110010000;
filter5[3][107] = 35'b11111110111101111000001111011010000;
filter5[3][108] = 35'b00000000011001010000111101111111100;
filter5[3][109] = 35'b11111011011101010100110010111000000;
filter5[3][110] = 35'b11111100111000011010011011101000000;
filter5[3][111] = 35'b11111111010101100111011111001101000;
filter5[3][112] = 35'b11111110101110001101001111000000000;
filter5[3][113] = 35'b00000000101000100111010001100110000;
filter5[3][114] = 35'b11111111101001010010001111010111100;
filter5[3][115] = 35'b00000000000001000111101111110010000;
filter5[3][116] = 35'b11111111100000011111001011010111000;
filter5[3][117] = 35'b00000010001000100010101000100100000;
filter5[3][118] = 35'b11111110001000101111111110111100000;
filter5[3][119] = 35'b11111111111100001001001010110000000;
filter5[3][120] = 35'b11111101001011101101000100101000000;
filter5[3][121] = 35'b00000010001010110010011110001000000;
filter5[3][122] = 35'b00000101010001100011111000101000000;
filter5[3][123] = 35'b00000101010001011101100110110000000;
filter5[3][124] = 35'b11111100010000100010101000001000000;
filter5[3][125] = 35'b11111101001011110001000001001100000;
filter5[3][126] = 35'b11111111011011111011111011001010000;
filter5[3][127] = 35'b11111010110111010010001101010000000;
filter5[3][128] = 35'b11111100001101101110011100101000000;
filter5[3][129] = 35'b11111000100011010010001111111000000;
filter5[3][130] = 35'b00000011010100101101010100001000000;
filter5[3][131] = 35'b00001000110101100000001000010000000;
filter5[3][132] = 35'b00000101100011010100110100010000000;
filter5[3][133] = 35'b00000110010100100101111100001000000;
filter5[3][134] = 35'b11101111010100111110001111000000000;
filter5[3][135] = 35'b11111000101001100111111010001000000;
filter5[3][136] = 35'b11110111101100111101110010100000000;
filter5[3][137] = 35'b00000110110100001011010011001000000;
filter5[3][138] = 35'b00000101010010111111111111001000000;
filter5[3][139] = 35'b11111011100111100000010110100000000;
filter5[3][140] = 35'b00000000000100110001110000101110111;
filter5[3][141] = 35'b00000001100110110101111011101010000;
filter5[3][142] = 35'b11111111100111100000111011011010000;
filter5[3][143] = 35'b11110101001110010011111001010000000;
filter5[3][144] = 35'b11111111001010010011011001110111000;
filter5[3][145] = 35'b11111111110110010010011110110110000;
filter5[3][146] = 35'b00000000101011110011110011110000000;
filter5[3][147] = 35'b00000010100011100110011100100000000;
filter5[3][148] = 35'b00000000011110001110110110101110000;
filter5[3][149] = 35'b11111111111101100011100011100010100;
filter5[3][150] = 35'b11111111100100000010010001000100100;
filter5[3][151] = 35'b11111101010101110000111000110100000;
filter5[3][152] = 35'b11111101111001001111110010100100000;
filter5[3][153] = 35'b11111110111010111001000000110010000;
filter5[3][154] = 35'b11111011111100011011000110111000000;
filter5[3][155] = 35'b00000011001011101111011101101100000;
filter5[3][156] = 35'b00000010010101101111010011110000000;
filter5[3][157] = 35'b00000010001010111010111010110100000;
filter5[3][158] = 35'b11111111001111100100011010000110000;
filter5[3][159] = 35'b11111011001010000110011110010000000;
filter5[3][160] = 35'b11111010101110100101000000001000000;
filter5[3][161] = 35'b11111100011101100101111000110000000;
filter5[3][162] = 35'b11111000001100001101101101010000000;
filter5[3][163] = 35'b00000111100011101111001011111000000;
filter5[3][164] = 35'b00000000001010111111001001111010100;
filter5[3][165] = 35'b11111111101100101110000000010001000;
filter5[3][166] = 35'b11110001011010011000110110110000000;
filter5[3][167] = 35'b11110110000010101000111001010000000;
filter5[3][168] = 35'b00000100110101101010011111010000000;
filter5[3][169] = 35'b11111000100111000001100000010000000;
filter5[3][170] = 35'b00000100000111010101001101111000000;
filter5[3][171] = 35'b11111110100101101010111100010000000;
filter5[3][172] = 35'b11111100000000100101001100100100000;
filter5[3][173] = 35'b11111001100110110111000101011000000;
filter5[3][174] = 35'b11101100100010110000110011100000000;
filter5[3][175] = 35'b11111010111111001001010011101000000;
filter5[3][176] = 35'b11101101010101100100000000100000000;
filter5[3][177] = 35'b00000011001000111111000010101100000;
filter5[3][178] = 35'b00000000100000001111100000011001000;
filter5[3][179] = 35'b11111101010000100011101111110000000;
filter5[3][180] = 35'b11111000110101110110101010010000000;
filter5[3][181] = 35'b11110111011011001110110101110000000;
filter5[3][182] = 35'b11110111011011110000100011000000000;
filter5[3][183] = 35'b00000000111100110101100110111110000;
filter5[3][184] = 35'b00000101011001110001100101110000000;
filter5[3][185] = 35'b00000110010010011111110011010000000;
filter5[3][186] = 35'b11110110101101000010100000000000000;
filter5[3][187] = 35'b00000111001010001011101001110000000;
filter5[3][188] = 35'b00000010001110001010010001010100000;
filter5[3][189] = 35'b11111010100111011010001111111000000;
filter5[3][190] = 35'b00001011101010100000011000100000000;
filter5[3][191] = 35'b11110101001010010000111111000000000;
filter5[3][192] = 35'b00000001011010011001110000110110000;
filter5[3][193] = 35'b11111011001001111111110001100000000;
filter5[3][194] = 35'b11111110100101000010100111110000000;
filter5[3][195] = 35'b00000001010011011101000111110010000;
filter5[3][196] = 35'b00000110010111011001110000001000000;
filter5[3][197] = 35'b00000101011001001001101010001000000;
filter5[3][198] = 35'b11110111010010001100110101100000000;
filter5[3][199] = 35'b11111001100011001111001000111000000;
filter5[3][200] = 35'b00000011000010110101001010111000000;
filter5[3][201] = 35'b11110011110011100110000011010000000;
filter5[3][202] = 35'b00000011101111101001111000101000000;
filter5[3][203] = 35'b00001010001100000110001100100000000;
filter5[3][204] = 35'b00000110100111110110000100111000000;
filter5[3][205] = 35'b00000001111011110101010010001010000;
filter5[3][206] = 35'b00000100110101100011000110110000000;
filter5[3][207] = 35'b11111111101110100110000100110110000;
filter5[3][208] = 35'b11111000000101000001110110000000000;
filter5[3][209] = 35'b11111101110011111110111011100100000;
filter5[3][210] = 35'b00000100011001111100000010110000000;
filter5[3][211] = 35'b00000010000001110001111011001100000;
filter5[3][212] = 35'b00000000011111001111100000110001000;
filter5[3][213] = 35'b11111100100000000101111100010100000;
filter5[3][214] = 35'b11111100110110011110000000110000000;
filter5[3][215] = 35'b11111110000100101010101010110000000;
filter5[3][216] = 35'b11111110100000101001000101001110000;
filter5[3][217] = 35'b11111100101100010100110011001000000;
filter5[3][218] = 35'b00000000101000110100110001000000000;
filter5[3][219] = 35'b00000011000011001011101011000100000;
filter5[3][220] = 35'b11111111100010011001100011101011100;
filter5[3][221] = 35'b11111111111100001110011100101000101;
filter5[3][222] = 35'b11111101011110111001110011001000000;
filter5[3][223] = 35'b11111011000001111101111011010000000;
filter5[3][224] = 35'b11111101001000110111101001111100000;
filter5[3][225] = 35'b00000010110101001010111010000100000;
filter5[3][226] = 35'b11111111000111001111111100110101000;
filter5[3][227] = 35'b11111111011000101010101100010011000;
filter5[3][228] = 35'b11111111010001100001001010100011000;
filter5[3][229] = 35'b00000100000100100001011000100000000;
filter5[3][230] = 35'b11111100011100000010111100000100000;
filter5[3][231] = 35'b11111011011000011011100101000000000;
filter5[3][232] = 35'b11111110010101001100110100101000000;
filter5[3][233] = 35'b00000010001111001111110111101100000;
filter5[3][234] = 35'b11111111101100100101101110101101100;
filter5[3][235] = 35'b00000000100001010110010001101111000;
filter5[3][236] = 35'b00000001001001101101100011101100000;
filter5[3][237] = 35'b11111101101001101110001110101000000;
filter5[3][238] = 35'b11111011110111000110110010100000000;
filter5[3][239] = 35'b11111010010110000010010001101000000;
filter5[3][240] = 35'b11111110010010001100100000000000000;
filter5[3][241] = 35'b00000001000001010100111110001110000;
filter5[3][242] = 35'b00000001100000100101100010110110000;
filter5[3][243] = 35'b11111111110001010111011010101010100;
filter5[3][244] = 35'b11111110011011010011000001011000000;
filter5[3][245] = 35'b11111111001110001111111110101011000;
filter5[3][246] = 35'b11111101110011111101101111100000000;
filter5[3][247] = 35'b11111011110000000000111111101000000;
filter5[3][248] = 35'b11111101101111110000001100011000000;
filter5[3][249] = 35'b00000011011110011010111110101000000;
filter5[3][250] = 35'b11111110001001011100001011100100000;
filter5[3][251] = 35'b11111111111010010100010001010010001;
filter5[3][252] = 35'b00000011100010001110110010001100000;
filter5[3][253] = 35'b00000000101111101010111001010101000;
filter5[3][254] = 35'b11111111001111101011001001110101000;
filter5[3][255] = 35'b00000010011101111011000011110000000;
filter5[3][256] = 35'b11111111001001101100111010111101000;
filter5[3][257] = 35'b11111101101100110101001001101000000;
filter5[3][258] = 35'b11111011001100011100111000111000000;
filter5[3][259] = 35'b00000011010111001001010110100100000;
filter5[3][260] = 35'b00000111110011010110001111010000000;
filter5[3][261] = 35'b11111011100000101100101101001000000;
filter5[3][262] = 35'b11111001010101011011111111110000000;
filter5[3][263] = 35'b00000000000011010000100011000000010;
filter5[3][264] = 35'b11111011101101111111111000010000000;
filter5[3][265] = 35'b11110110101100100101001100110000000;
filter5[3][266] = 35'b00000001000011110001101000001110000;
filter5[3][267] = 35'b00000101110100000100010010100000000;
filter5[3][268] = 35'b11111111100001110100010101000001000;
filter5[3][269] = 35'b11111111110101001011101110110011100;
filter5[3][270] = 35'b11110111000001101010101110110000000;
filter5[3][271] = 35'b11111101001101100110010100011000000;
filter5[3][272] = 35'b11111110000101111010000101010000000;
filter5[3][273] = 35'b11111111110111011010001111101011010;
filter5[3][274] = 35'b00000010101100010101101111010100000;
filter5[3][275] = 35'b00000000100010000101001101111100000;
filter5[3][276] = 35'b11111110011010101111100010100010000;
filter5[3][277] = 35'b00000000010111110000101000011011000;
filter5[3][278] = 35'b00000000100011100010000010001010000;
filter5[3][279] = 35'b11111001011011111101011011000000000;
filter5[3][280] = 35'b00000001001101111011101011110000000;
filter5[3][281] = 35'b00000000110011110000100000111010000;
filter5[3][282] = 35'b00000001100111000101001110100110000;
filter5[3][283] = 35'b11111110000110100011000000000010000;
filter5[3][284] = 35'b11111110100001000110110000100100000;
filter5[3][285] = 35'b00000000101111110001001110110110000;
filter5[3][286] = 35'b00000000001001110101001100000011000;
filter5[3][287] = 35'b11111101000100011000000111100000000;
filter5[3][288] = 35'b11111111001110100111001111100111000;
filter5[3][289] = 35'b00000010000101001000101010101000000;
filter5[3][290] = 35'b00000000001000011000010101010001000;
filter5[3][291] = 35'b00000011011010001101101100110100000;
filter5[3][292] = 35'b11111111100011010110111111100110100;
filter5[3][293] = 35'b11111110010100110101110001001010000;
filter5[3][294] = 35'b00000001000011110101000000011010000;
filter5[3][295] = 35'b11111110111110111011010011110100000;
filter5[3][296] = 35'b11111101011011010110011100111100000;
filter5[3][297] = 35'b00000001010100111000000100000010000;
filter5[3][298] = 35'b11111100111001111110111000101000000;
filter5[3][299] = 35'b00000100110110111111101001111000000;
filter5[3][300] = 35'b11111110111100101101110001000100000;
filter5[3][301] = 35'b11111110001011011111001011101100000;
filter5[3][302] = 35'b00000001010001010011100010100110000;
filter5[3][303] = 35'b00000001110001111100011110000100000;
filter5[3][304] = 35'b11111110101001011001011110111000000;
filter5[3][305] = 35'b00000001101110110011000001101010000;
filter5[3][306] = 35'b00000010000110100110100010000000000;
filter5[3][307] = 35'b00000010000110011100110110001000000;
filter5[3][308] = 35'b11111110011100011010110110001000000;
filter5[3][309] = 35'b00000001001010010110101100010110000;
filter5[3][310] = 35'b11111110000001000101000110110010000;
filter5[3][311] = 35'b00000010001000100111010001001000000;
filter5[3][312] = 35'b11111011010001000010100001111000000;
filter5[3][313] = 35'b00000110010001000111011111001000000;
filter5[3][314] = 35'b00000011110110111101100010001100000;
filter5[3][315] = 35'b11111100110101000001010101010100000;
filter5[3][316] = 35'b11111101001000011000101110101100000;
filter5[3][317] = 35'b11111100000100010110111011011100000;
filter5[3][318] = 35'b00000000000000000010101010100101110;
filter5[3][319] = 35'b11111010011011000001110100001000000;
filter5[3][320] = 35'b11111000010000000110111010100000000;
filter5[3][321] = 35'b11111110001110110110111000110000000;
filter5[3][322] = 35'b00000110000011011000100010101000000;
filter5[3][323] = 35'b00000111000011110101100110100000000;
filter5[3][324] = 35'b00000011010011100101000010110000000;
filter5[3][325] = 35'b00000100011000101001011111110000000;
filter5[3][326] = 35'b11110111011001111001110000110000000;
filter5[3][327] = 35'b11111011101110000011111010001000000;
filter5[3][328] = 35'b00000011011000110010101000101000000;
filter5[3][329] = 35'b00000100010100010100110110010000000;
filter5[3][330] = 35'b00000011000011010001001111101100000;
filter5[3][331] = 35'b00000011011000101010001001110100000;
filter5[3][332] = 35'b00000011010001110110111011001100000;
filter5[3][333] = 35'b00000010011110011110010101100000000;
filter5[3][334] = 35'b11111111111001001111111111111000010;
filter5[3][335] = 35'b11111101011111001010011010111100000;
filter5[3][336] = 35'b11111110010011110000011010111100000;
filter5[3][337] = 35'b00000001011100010000111010010110000;
filter5[3][338] = 35'b00000011011001000101000000101000000;
filter5[3][339] = 35'b11111100100001001000000111110000000;
filter5[3][340] = 35'b11111110001001010101101011110010000;
filter5[3][341] = 35'b11111101110000100000000111010100000;
filter5[3][342] = 35'b11111101111010000011010101101100000;
filter5[3][343] = 35'b11111111001111010101110110100110000;
filter5[3][344] = 35'b00000000101001111100100100010000000;
filter5[3][345] = 35'b00000100101100000100011000101000000;
filter5[3][346] = 35'b00000001111011001111001000100100000;
filter5[3][347] = 35'b11111100001111000100101001001100000;
filter5[3][348] = 35'b11111100111000101000111111101100000;
filter5[3][349] = 35'b11111101101100010010010101011000000;
filter5[3][350] = 35'b11111110001111100010011111010110000;
filter5[3][351] = 35'b11111110110101100111100101001100000;
filter5[3][352] = 35'b00000010100010101011000111101000000;
filter5[3][353] = 35'b00000101100110101110011110010000000;
filter5[3][354] = 35'b11111011011101010010010100000000000;
filter5[3][355] = 35'b00000000011100111001110011110001000;
filter5[3][356] = 35'b11111111011011111101001111011100000;
filter5[3][357] = 35'b00000101000110100110001110110000000;
filter5[3][358] = 35'b11111010001110011011100001100000000;
filter5[3][359] = 35'b11111111101011100011000101111000100;
filter5[3][360] = 35'b00000001001111111110000110100100000;
filter5[3][361] = 35'b00000010000101010111100010110100000;
filter5[3][362] = 35'b11111111000101110101011110101111000;
filter5[3][363] = 35'b11111101000010001111100011110000000;
filter5[3][364] = 35'b00000001011000110101011110101010000;
filter5[3][365] = 35'b11111101101000100111010101111000000;
filter5[3][366] = 35'b11111100101001011100001101001000000;
filter5[3][367] = 35'b11111101101001000100101010100000000;
filter5[3][368] = 35'b00000000111000000011011011101011000;
filter5[3][369] = 35'b11111100101000110101111011011000000;
filter5[3][370] = 35'b00000000100000110010110111000101000;
filter5[3][371] = 35'b00000000011111110100011110010011000;
filter5[3][372] = 35'b00000011101101001010100101001100000;
filter5[3][373] = 35'b11111110000111001111000110101100000;
filter5[3][374] = 35'b11111100011101110100110010011100000;
filter5[3][375] = 35'b11111100101101011110011010110000000;
filter5[3][376] = 35'b00000011001000011001101111001100000;
filter5[3][377] = 35'b00000001001110011001111110000010000;
filter5[3][378] = 35'b11111111111010110011001000111010010;
filter5[3][379] = 35'b00000010101011010000100110100100000;
filter5[3][380] = 35'b00000001011111000111100111001000000;
filter5[3][381] = 35'b00000001010011110001110000111110000;
filter5[3][382] = 35'b00000010000100110100011011001000000;
filter5[3][383] = 35'b00000010000101001111101101010000000;
filter5[3][384] = 35'b11111101010000001010000111011100000;
filter5[3][385] = 35'b11111100010010011011000110101100000;
filter5[3][386] = 35'b00000001100000011101111011100110000;
filter5[3][387] = 35'b00000000110000111100001000011101000;
filter5[3][388] = 35'b00000010000011011010000010001000000;
filter5[3][389] = 35'b11111110000110000011000001011000000;
filter5[3][390] = 35'b00000011101000010001010001110100000;
filter5[3][391] = 35'b11111101011111001110010110010000000;
filter5[3][392] = 35'b00000011110011111011000001011100000;
filter5[3][393] = 35'b00000010010010100111100111100000000;
filter5[3][394] = 35'b00000010100010100000100101010000000;
filter5[3][395] = 35'b11111101001000000100001110011000000;
filter5[3][396] = 35'b11111111000111011011101000111100000;
filter5[3][397] = 35'b00000010110000001011111000101100000;
filter5[3][398] = 35'b00000001110111010110001000110010000;
filter5[3][399] = 35'b00000100110011000000000111100000000;
filter5[3][400] = 35'b00000000101100001000111110010011000;
filter5[3][401] = 35'b00000010101101111000011101001100000;
filter5[3][402] = 35'b00000000001010010101001111010110100;
filter5[3][403] = 35'b00000001100101110000101101011000000;
filter5[3][404] = 35'b11111100110100010001111110000000000;
filter5[3][405] = 35'b11111111111000110111011111111010010;
filter5[3][406] = 35'b00000000110100101010111011101001000;
filter5[3][407] = 35'b00000010111100101100110010001000000;
filter5[3][408] = 35'b11111110101000110011011110000100000;
filter5[3][409] = 35'b00000000000011101010001001011110111;
filter5[3][410] = 35'b11111101101110001001111111111100000;
filter5[3][411] = 35'b11111001101100100110110101101000000;
filter5[3][412] = 35'b00000001001100001100111100100010000;
filter5[3][413] = 35'b11111111101001111110010101001011000;
filter5[3][414] = 35'b00000011111001100010001111101100000;
filter5[3][415] = 35'b11111111101100101110000000001100100;
filter5[3][416] = 35'b00000000111000010111101100101011000;
filter5[3][417] = 35'b00000010010110110000111000110000000;
filter5[3][418] = 35'b00000001110101001100111111101110000;
filter5[3][419] = 35'b11111011010011111001101001010000000;
filter5[3][420] = 35'b11111111010101011000000101010110000;
filter5[3][421] = 35'b11111011001101101010100011010000000;
filter5[3][422] = 35'b00000011111000001001111110110000000;
filter5[3][423] = 35'b11111111110111110010010111001110100;
filter5[3][424] = 35'b00000001010101110111000101000110000;
filter5[3][425] = 35'b11111011011010100100111001001000000;
filter5[3][426] = 35'b11111101010111110001101001100100000;
filter5[3][427] = 35'b11111011010110001101010111100000000;
filter5[3][428] = 35'b11111101000010100011001110111000000;
filter5[3][429] = 35'b00000010100000001100000011101000000;
filter5[3][430] = 35'b11111111011001111001001010000001000;
filter5[3][431] = 35'b00000010000110000010101110011000000;
filter5[3][432] = 35'b00000000111010110101001000110100000;
filter5[3][433] = 35'b00000001010000010011111010101000000;
filter5[3][434] = 35'b00000000001001010000110011000010010;
filter5[3][435] = 35'b11111101001111111001101010000100000;
filter5[3][436] = 35'b00000001111010011000001000011010000;
filter5[3][437] = 35'b11111110001111010000000010000110000;
filter5[3][438] = 35'b11111111000111010001011100000010000;
filter5[3][439] = 35'b00000010010000111100001001011100000;
filter5[3][440] = 35'b11111011011000000000010011100000000;
filter5[3][441] = 35'b00000100101000100010010111010000000;
filter5[3][442] = 35'b11111110100010111000000010000010000;
filter5[3][443] = 35'b00000010101010001110110000101000000;
filter5[3][444] = 35'b00000001110010100000000111111100000;
filter5[3][445] = 35'b11111111110011000101101001101101010;
filter5[3][446] = 35'b00000010001100001100011011100000000;
filter5[3][447] = 35'b11111111000000001000011011110010000;
filter5[3][448] = 35'b00000010000101100101101000110000000;
filter5[3][449] = 35'b00000001001011101100110110000110000;
filter5[3][450] = 35'b00000010000100011111000001011100000;
filter5[3][451] = 35'b11111001111100110001011110111000000;
filter5[3][452] = 35'b11111100010011101110001101010000000;
filter5[3][453] = 35'b00000000100000101010010011111100000;
filter5[3][454] = 35'b00000100101000110011010111110000000;
filter5[3][455] = 35'b00000010111111001100101111010100000;
filter5[3][456] = 35'b11111110110111100110011001010110000;
filter5[3][457] = 35'b11111101010000000011000101101100000;
filter5[3][458] = 35'b11111101110110111011100111111100000;
filter5[3][459] = 35'b11111011001000111000010001110000000;
filter5[3][460] = 35'b11111001010101101011000100100000000;
filter5[3][461] = 35'b11111001011111001001011010110000000;
filter5[3][462] = 35'b11111011011000001101000100001000000;
filter5[3][463] = 35'b00000000001110000001100010001100010;
filter5[3][464] = 35'b11111110001000111010111100010000000;
filter5[3][465] = 35'b11110110010010011111100000110000000;
filter5[3][466] = 35'b11111100010011111000011111100000000;
filter5[3][467] = 35'b11111101000100011101101011110000000;
filter5[3][468] = 35'b11110111011110110101001011000000000;
filter5[3][469] = 35'b11110010011101100001010010000000000;
filter5[3][470] = 35'b11111100000010101000110100001100000;
filter5[3][471] = 35'b00000011000001111011100001110000000;
filter5[3][472] = 35'b11100110110101001000111011000000000;
filter5[3][473] = 35'b11101001011010001100001001000000000;
filter5[3][474] = 35'b11111110000101010001100111100010000;
filter5[3][475] = 35'b11111100111111000000111000111000000;
filter5[3][476] = 35'b00000011101001111010011101010000000;
filter5[3][477] = 35'b00000011000101010011111111101000000;
filter5[3][478] = 35'b00000000111010110001110011011010000;
filter5[3][479] = 35'b00000010101111101101110001001000000;
filter5[3][480] = 35'b11110100100111010100011000000000000;
filter5[3][481] = 35'b11101110101011110011010000000000000;
filter5[3][482] = 35'b11111000111000110110001001010000000;
filter5[3][483] = 35'b00000001010111111100011110010010000;
filter5[3][484] = 35'b00000000101001100011110001001010000;
filter5[3][485] = 35'b11111110101100101010101001000100000;
filter5[3][486] = 35'b00000010111010100110010000010000000;
filter5[3][487] = 35'b00000001101000010011010000111010000;
filter5[3][488] = 35'b00000101001000011100011101110000000;
filter5[3][489] = 35'b11111111011000011111000010110111000;
filter5[3][490] = 35'b11111111011100010000100110000100000;
filter5[3][491] = 35'b11111100000000101111001000000100000;
filter5[3][492] = 35'b11111101111101110110000111101100000;
filter5[3][493] = 35'b11111101001011100101010110010100000;
filter5[3][494] = 35'b00000001000000101010000000101100000;
filter5[3][495] = 35'b11111111110110001111010111101100100;
filter5[3][496] = 35'b00000010001000000101010001101000000;
filter5[3][497] = 35'b00000100001110000001110001110000000;
filter5[3][498] = 35'b00000000101011111100000100001001000;
filter5[3][499] = 35'b11111100011011000100100001001100000;
filter5[3][500] = 35'b11111110110110010000011000101100000;
filter5[3][501] = 35'b11110111101101000111010011100000000;
filter5[3][502] = 35'b00000001010111111011111100100110000;
filter5[3][503] = 35'b00000000100000011111100110001100000;
filter5[3][504] = 35'b00000100001001011101010000011000000;
filter5[3][505] = 35'b11111111110010101010000011001010100;
filter5[3][506] = 35'b00000010000100111100010111100000000;
filter5[3][507] = 35'b00000001011101001101011101110110000;
filter5[3][508] = 35'b00000010001010001101100101111100000;
filter5[3][509] = 35'b11111111001101010111101101011010000;
filter5[3][510] = 35'b00000001111010101100111010001100000;
filter5[3][511] = 35'b11111110101001001110001110001000000;
filter5[3][512] = 35'b00000000101000010010111010101100000;
filter5[3][513] = 35'b11111111101110110001001110001111000;
filter5[3][514] = 35'b00000001100100001111100101110010000;
filter5[3][515] = 35'b00000010100111000000101001000100000;
filter5[3][516] = 35'b11111111001100100111100101001010000;
filter5[3][517] = 35'b00000000111110010011110110100100000;
filter5[3][518] = 35'b00000000100110011110101001000111000;
filter5[3][519] = 35'b11111000101111111010110110111000000;
filter5[3][520] = 35'b00000010101111100110001101100000000;
filter5[3][521] = 35'b00000010010011100100111000010000000;
filter5[3][522] = 35'b11111110110000001101111011101010000;
filter5[3][523] = 35'b00000000100011011101000110011010000;
filter5[3][524] = 35'b00000000010111101011100011001100100;
filter5[3][525] = 35'b00000000110010101110111101111000000;
filter5[3][526] = 35'b11111111001100110101001001000111000;
filter5[3][527] = 35'b00000001100010100100110110110110000;
filter5[3][528] = 35'b11111010011010111110000011100000000;
filter5[3][529] = 35'b11111111110101110111110100010010010;
filter5[3][530] = 35'b00000100111000011101001101110000000;
filter5[3][531] = 35'b11111101110101101110110111000000000;
filter5[3][532] = 35'b00000000010001011000010011110110100;
filter5[3][533] = 35'b00000001101001010001100011011000000;
filter5[3][534] = 35'b00000100111100010000101001001000000;
filter5[3][535] = 35'b11111110110100010111110100000010000;
filter5[3][536] = 35'b11111110011100110100001010000100000;
filter5[3][537] = 35'b00000100001001000000101000101000000;
filter5[3][538] = 35'b11111111111110100000011010111011100;
filter5[3][539] = 35'b11111110000111111011001101010010000;
filter5[3][540] = 35'b11111011101100110010111001110000000;
filter5[3][541] = 35'b11111111000001000001100010100100000;
filter5[3][542] = 35'b11111110101001010010000011111000000;
filter5[3][543] = 35'b11111111011010110101100010101000000;
filter5[3][544] = 35'b11111100000101101101001000110100000;
filter5[3][545] = 35'b00000001000010110111010000111000000;
filter5[3][546] = 35'b00000001011111000010101011101010000;
filter5[3][547] = 35'b11111110101101010000011010010110000;
filter5[3][548] = 35'b11111110011010101000101101011010000;
filter5[3][549] = 35'b00000000001010001101000111111100100;
filter5[3][550] = 35'b11111110011000011111101000000000000;
filter5[3][551] = 35'b00000011110011000111111011011000000;
filter5[3][552] = 35'b11111101110100010110000000010000000;
filter5[3][553] = 35'b00000010110100001100010010010100000;
filter5[3][554] = 35'b11111000010011110100010000101000000;
filter5[3][555] = 35'b00000000100001100001001011001000000;
filter5[3][556] = 35'b00000000110000011100001000100011000;
filter5[3][557] = 35'b11111111001110001100111110101100000;
filter5[3][558] = 35'b11111100100001010000111101000100000;
filter5[3][559] = 35'b00000010111101110011101110110000000;
filter5[3][560] = 35'b00000100101100011101001110010000000;
filter5[3][561] = 35'b11111110110011010100100010000100000;
filter5[3][562] = 35'b00000001011001100111101011111000000;
filter5[3][563] = 35'b11111111110001010101110111010110100;
filter5[3][564] = 35'b00000100111000111010100000010000000;
filter5[3][565] = 35'b11111101111110010100100011011100000;
filter5[3][566] = 35'b11111111001011101000100100001000000;
filter5[3][567] = 35'b00000010001001111011110001010000000;
filter5[3][568] = 35'b11111101110101011011011011011100000;
filter5[3][569] = 35'b11111110001011000000010000010010000;
filter5[3][570] = 35'b00000011000110010010010011101000000;
filter5[3][571] = 35'b00000001101100000010011000011110000;
filter5[3][572] = 35'b00000001100000000000101100100110000;
filter5[3][573] = 35'b00000000110011110100001000101100000;
filter5[3][574] = 35'b00000011011010101010010110111000000;
filter5[3][575] = 35'b00000001111011101001101100001110000;
filter5[3][576] = 35'b11111101001111010010101001101100000;
filter5[3][577] = 35'b00000000000011110001001010000010100;
filter5[3][578] = 35'b00000100000010101000100110011000000;
filter5[3][579] = 35'b00000000101010001001100101001010000;
filter5[3][580] = 35'b00000001100111101001010011110110000;
filter5[3][581] = 35'b00000100011001010001101100100000000;
filter5[3][582] = 35'b00000110001000100100100010011000000;
filter5[3][583] = 35'b11111100010001000001000100111100000;
filter5[3][584] = 35'b00000001000001000000011011101010000;
filter5[3][585] = 35'b11111000111011010101000000110000000;
filter5[3][586] = 35'b00000000011100010101010011001011100;
filter5[3][587] = 35'b00000100001101111011100111101000000;
filter5[3][588] = 35'b00000001100101010101010001111010000;
filter5[3][589] = 35'b00000100110110011000100011100000000;
filter5[3][590] = 35'b00000001100110100100000000111100000;
filter5[3][591] = 35'b00000101011100101100011010111000000;
filter5[3][592] = 35'b11111011100001111101010010111000000;
filter5[3][593] = 35'b00000000001101001111110001010100010;
filter5[3][594] = 35'b11111111010010101110100011100111000;
filter5[3][595] = 35'b00000000111110110010100001001011000;
filter5[3][596] = 35'b11111110101101010001010011110010000;
filter5[3][597] = 35'b11111101111001011100010101111000000;
filter5[3][598] = 35'b11111111101000100111011110100111100;
filter5[3][599] = 35'b11111111100011001000000001100110100;
filter5[3][600] = 35'b11111100100000101100011001100000000;
filter5[3][601] = 35'b11111101010100111110100001000000000;
filter5[3][602] = 35'b11111110111110011001001000001110000;
filter5[3][603] = 35'b11111110110101010001000011101000000;
filter5[3][604] = 35'b11111111110101001100101001101110100;
filter5[3][605] = 35'b11111111111101010101011100000011000;
filter5[3][606] = 35'b11111111111010110110000010001100000;
filter5[3][607] = 35'b11111011010010000010011101011000000;
filter5[3][608] = 35'b11110010100101010010010100100000000;
filter5[3][609] = 35'b00000001010110110110110000100000000;
filter5[3][610] = 35'b00000001010001010111001100011100000;
filter5[3][611] = 35'b00000011001110101001011100111100000;
filter5[3][612] = 35'b00000000000110010110010010100110010;
filter5[3][613] = 35'b00000011011101000011010001010000000;
filter5[3][614] = 35'b11111110010001000000111111110100000;
filter5[3][615] = 35'b00000000011010111000100100100001100;
filter5[3][616] = 35'b11111001010100001111001010111000000;
filter5[3][617] = 35'b11111101111110110011010000101000000;
filter5[3][618] = 35'b00000010001111011001110001110100000;
filter5[3][619] = 35'b00000001001101101110111010011100000;
filter5[3][620] = 35'b00000000101111111010001000111010000;
filter5[3][621] = 35'b11111110110001110001111011010010000;
filter5[3][622] = 35'b11111011011100001011000001101000000;
filter5[3][623] = 35'b11111110110111101011111111101000000;
filter5[3][624] = 35'b11111110011011001100110010011000000;
filter5[3][625] = 35'b00000000011010101111101100110100000;
filter5[3][626] = 35'b00000011001011010001010001101000000;
filter5[3][627] = 35'b00000001100000001110111001110110000;
filter5[3][628] = 35'b00000000010010011000111110000000000;
filter5[3][629] = 35'b11111110111000111000010011101000000;
filter5[3][630] = 35'b00000000001100100110001111011011010;
filter5[3][631] = 35'b00000000011010001101000001101110100;
filter5[3][632] = 35'b11111111110010101111001011000011100;
filter5[3][633] = 35'b11111101110100010111100001111100000;
filter5[3][634] = 35'b00000001001110011111011110000110000;
filter5[3][635] = 35'b11111101110010110111111011100000000;
filter5[3][636] = 35'b00000001100000100000000010000000000;
filter5[3][637] = 35'b11111101110011111110100011000100000;
filter5[3][638] = 35'b00000001101111111001111100110010000;
filter5[3][639] = 35'b11111110011100010110110010101110000;
filter5[3][640] = 35'b00000000011000101100011100101011100;
filter5[3][641] = 35'b11111100111101110011011011011100000;
filter5[3][642] = 35'b11111011001100011010011111000000000;
filter5[3][643] = 35'b11110110110010011010110011100000000;
filter5[3][644] = 35'b11111101100101111111110101001000000;
filter5[3][645] = 35'b00000100101011100010100110100000000;
filter5[3][646] = 35'b11111101010011100000101101111000000;
filter5[3][647] = 35'b11110100011001101011111101010000000;
filter5[3][648] = 35'b00000001000111110010101001011110000;
filter5[3][649] = 35'b11111010001010010001110010111000000;
filter5[3][650] = 35'b11111101000000101110111101011100000;
filter5[3][651] = 35'b00000000100011001000111100110100000;
filter5[3][652] = 35'b00000001010100110011000111011110000;
filter5[3][653] = 35'b00000001111101101100100010110000000;
filter5[3][654] = 35'b00000000001011011011011001011111100;
filter5[3][655] = 35'b11111011101000111011110110111000000;
filter5[3][656] = 35'b00000001100011111010100011001110000;
filter5[3][657] = 35'b00000100001011111100110010010000000;
filter5[3][658] = 35'b00000101000100010100010010100000000;
filter5[3][659] = 35'b11111110100110101011001110001100000;
filter5[3][660] = 35'b11111101011111011000010001010100000;
filter5[3][661] = 35'b11111101010010000000101000011000000;
filter5[3][662] = 35'b00000100110011100101011011111000000;
filter5[3][663] = 35'b11111110110010010001110100110100000;
filter5[3][664] = 35'b00000101101011001100101101111000000;
filter5[3][665] = 35'b00000000001010110001111110101001100;
filter5[3][666] = 35'b11111111001100100111000010010011000;
filter5[3][667] = 35'b11111111100011110000100001010111100;
filter5[3][668] = 35'b00000000001000110111011001110010110;
filter5[3][669] = 35'b00000000000101011100101011101100101;
filter5[3][670] = 35'b11111111101111000110110011100111100;
filter5[3][671] = 35'b00000000100000001101010101000010000;
filter5[3][672] = 35'b11111101011000101100101101010000000;
filter5[3][673] = 35'b00000101000101000001111000011000000;
filter5[3][674] = 35'b11111001100000001001100101001000000;
filter5[3][675] = 35'b00000000000011100111111100111101000;
filter5[3][676] = 35'b11111110001010010000010110000000000;
filter5[3][677] = 35'b11111111000010111101101101001000000;
filter5[3][678] = 35'b00000001101111111111000100100010000;
filter5[3][679] = 35'b00000001001010010000110111101000000;
filter5[3][680] = 35'b00000111011110100010100100110000000;
filter5[3][681] = 35'b00000000111000100101001010101011000;
filter5[3][682] = 35'b11111001101101111110110110100000000;
filter5[3][683] = 35'b11111110110110010100011111101110000;
filter5[3][684] = 35'b11111110110011000100101101010000000;
filter5[3][685] = 35'b00000010010001100001111100110000000;
filter5[3][686] = 35'b11111110111011100101011110001100000;
filter5[3][687] = 35'b00000010110011010100110101011000000;
filter5[3][688] = 35'b11111111101010101110011111111101000;
filter5[3][689] = 35'b00000010011100111001001010010000000;
filter5[3][690] = 35'b11111111110111001111001101000011100;
filter5[3][691] = 35'b11111110010111011010111000011000000;
filter5[3][692] = 35'b11111100101110101001000000101000000;
filter5[3][693] = 35'b11111110110100000010101100011100000;
filter5[3][694] = 35'b00000010000110101000110101011100000;
filter5[3][695] = 35'b00000010010100000100001011010100000;
filter5[3][696] = 35'b11111111110010011000101110101010000;
filter5[3][697] = 35'b00000001011010010011001010101000000;
filter5[3][698] = 35'b00000000001100111010010011101010000;
filter5[3][699] = 35'b00000000111100011111110010000111000;
filter5[3][700] = 35'b00000010110110010111010101011000000;
filter5[3][701] = 35'b11111111001000011111000010110010000;
filter5[3][702] = 35'b00000100011011010101111101111000000;
filter5[3][703] = 35'b11111111001011101010111011110001000;
filter5[3][704] = 35'b11111110010010000010110011010110000;
filter5[3][705] = 35'b11111110001100011011111001000100000;
filter5[3][706] = 35'b11111111011001111101001101101001000;
filter5[3][707] = 35'b00000010100011100111010000000000000;
filter5[3][708] = 35'b00000010000100110001100010001100000;
filter5[3][709] = 35'b11111111101101001111101101011010000;
filter5[3][710] = 35'b11111111010110101110110000111010000;
filter5[3][711] = 35'b11111111000000111001010010010001000;
filter5[3][712] = 35'b11111110000111100010100000011000000;
filter5[3][713] = 35'b00000000101010001010000110011001000;
filter5[3][714] = 35'b00000011001110000101011111001100000;
filter5[3][715] = 35'b11111101101001110001111011011000000;
filter5[3][716] = 35'b00000010100100101001000011010100000;
filter5[3][717] = 35'b11111101110011111000011101000100000;
filter5[3][718] = 35'b00000010001001101111111110010000000;
filter5[3][719] = 35'b11111111111110101110111010100011101;
filter5[3][720] = 35'b11111111000101011010010000000110000;
filter5[3][721] = 35'b11111011010000101100111101010000000;
filter5[3][722] = 35'b00000000001010011010100100010110010;
filter5[3][723] = 35'b11111110110101011111110000011100000;
filter5[3][724] = 35'b00000000001110110001111010110000010;
filter5[3][725] = 35'b11111010101001110101011100000000000;
filter5[3][726] = 35'b11111100111101110100100101111100000;
filter5[3][727] = 35'b11111111000010101110011100100010000;
filter5[3][728] = 35'b11111101101111110001010100001000000;
filter5[3][729] = 35'b11111110010111101101101011001010000;
filter5[3][730] = 35'b00000011001110110001010111110100000;
filter5[3][731] = 35'b00000100011001011000110100100000000;
filter5[3][732] = 35'b00000001000100111000101111111110000;
filter5[3][733] = 35'b11111110110111100001011011111010000;
filter5[3][734] = 35'b00000000111010100001011111000111000;
filter5[3][735] = 35'b11111101101010111001111011000100000;
filter5[3][736] = 35'b00000011000001001000101010000100000;
filter5[3][737] = 35'b00000010101100000111101011000000000;
filter5[3][738] = 35'b11111011100000000001111110101000000;
filter5[3][739] = 35'b00000000101100111000100000101010000;
filter5[3][740] = 35'b00000010100010000000000111010000000;
filter5[3][741] = 35'b11111100110111001110100110101000000;
filter5[3][742] = 35'b11111101100011010100110001011100000;
filter5[3][743] = 35'b11111110101111010110100000110000000;
filter5[3][744] = 35'b00000001100001010101000010101110000;
filter5[3][745] = 35'b00000011011100001011110110001100000;
filter5[3][746] = 35'b11111110010010100111101010000000000;
filter5[3][747] = 35'b11111110101010101011100000000010000;
filter5[3][748] = 35'b00000000001111010001111010000011100;
filter5[3][749] = 35'b00000001000110001111010000100100000;
filter5[3][750] = 35'b11111100001110111001101001010100000;
filter5[3][751] = 35'b11111111100000001011111011001100000;
filter5[3][752] = 35'b11111011100000111100100111100000000;
filter5[3][753] = 35'b00000100000100001011001000101000000;
filter5[3][754] = 35'b00000011001010011001000011000000000;
filter5[3][755] = 35'b11111110100011000001011101111110000;
filter5[3][756] = 35'b11111111010010110111100011001110000;
filter5[3][757] = 35'b00000000011101110100001010011001100;
filter5[3][758] = 35'b11111100110101010011001100000000000;
filter5[3][759] = 35'b11111011010101011001101100000000000;
filter5[3][760] = 35'b11111001100000011011101000101000000;
filter5[3][761] = 35'b00000001101111110011110111101110000;
filter5[3][762] = 35'b00000000001011011111101010111000110;
filter5[3][763] = 35'b00000011101100111110100110101100000;
filter5[3][764] = 35'b00000000001100100000110101100101010;
filter5[3][765] = 35'b11111110111111101010101111000010000;
filter5[3][766] = 35'b00000000110000000010111000111001000;
filter5[3][767] = 35'b11111101000010110001000111000000000;
filter5[3][768] = 35'b11111101001011011111011100011100000;
filter5[3][769] = 35'b00000001111001110100011110000000000;
filter5[3][770] = 35'b00000101110100100000001111110000000;
filter5[3][771] = 35'b00000010010010100111101101000000000;
filter5[3][772] = 35'b11111000111100001010000101011000000;
filter5[3][773] = 35'b00000010111001110010011001000100000;
filter5[3][774] = 35'b11111111110110111000001010101001100;
filter5[3][775] = 35'b11111110100100000111110111100010000;
filter5[3][776] = 35'b00000001111111101100110101010100000;
filter5[3][777] = 35'b00000110000110101001010011100000000;
filter5[3][778] = 35'b11111110011011010010111101101000000;
filter5[3][779] = 35'b00000000011101011011011110100100100;
filter5[3][780] = 35'b11111110001110011101010010000110000;
filter5[3][781] = 35'b11111001011000110101100100110000000;
filter5[3][782] = 35'b00000100100100101101101000010000000;
filter5[3][783] = 35'b00000001011000000001010001010100000;
filter5[3][784] = 35'b00000011100000110101000110000000000;
filter5[3][785] = 35'b00000110000000010001111001111000000;
filter5[3][786] = 35'b00000111111001000010101111111000000;
filter5[3][787] = 35'b11111100000100001001010111101000000;
filter5[3][788] = 35'b11111011101010010110101111000000000;
filter5[3][789] = 35'b11111011101001010010101010010000000;
filter5[3][790] = 35'b11111100011001101000100101111100000;
filter5[3][791] = 35'b00000010100100101010100011010100000;
filter5[3][792] = 35'b00000010010100011101010110101100000;
filter5[3][793] = 35'b00000101010101101101101011010000000;
filter5[3][794] = 35'b11111011110101001001011010000000000;
filter5[3][795] = 35'b11111111100110100011100001110011100;
filter5[3][796] = 35'b00000100001110110011100010110000000;
filter5[3][797] = 35'b00000101010100111000111100100000000;
filter5[3][798] = 35'b11111011000101001011011000010000000;
filter5[3][799] = 35'b00000110110010000011011110100000000;
filter5[3][800] = 35'b00000010000000101001101101011000000;
filter5[3][801] = 35'b11111100001000111100100110111000000;
filter5[3][802] = 35'b11111100110000011101111111110100000;
filter5[3][803] = 35'b11111001110011111001110100101000000;
filter5[3][804] = 35'b00000100100110111010100001000000000;
filter5[3][805] = 35'b00000010110001000101010011100100000;
filter5[3][806] = 35'b11111111000111011000100000000100000;
filter5[3][807] = 35'b00000010001111101111111100101100000;
filter5[3][808] = 35'b00000100001011001011001100100000000;
filter5[3][809] = 35'b11110101000011111010011001000000000;
filter5[3][810] = 35'b11111000010011010101001001110000000;
filter5[3][811] = 35'b11111100000111101110101101100100000;
filter5[3][812] = 35'b11111110001010000011100001101100000;
filter5[3][813] = 35'b11111101100110001100110101101100000;
filter5[3][814] = 35'b00000001000101001011011110101000000;
filter5[3][815] = 35'b11111110101100100110000000100100000;
filter5[3][816] = 35'b00000000101011011011101110001110000;
filter5[3][817] = 35'b11111100011010000111010010110100000;
filter5[3][818] = 35'b11111101100101110001100110100100000;
filter5[3][819] = 35'b11111111011111010110101011011111000;
filter5[3][820] = 35'b00000010110100010000000101101100000;
filter5[3][821] = 35'b11111001101011001011111011000000000;
filter5[3][822] = 35'b11111110001010011000100101010010000;
filter5[3][823] = 35'b00000011011101101110001000110000000;
filter5[3][824] = 35'b00000011100000110111101100100000000;
filter5[3][825] = 35'b00000011000001100001101111111100000;
filter5[3][826] = 35'b00000100101111111111100101010000000;
filter5[3][827] = 35'b00000000111111100111000101000011000;
filter5[3][828] = 35'b11111101111011010001100000101100000;
filter5[3][829] = 35'b11111111100001100010001000001100000;
filter5[3][830] = 35'b00000001010010100001000100111000000;
filter5[3][831] = 35'b00000000000111010110001010011110111;
filter5[3][832] = 35'b00000000000000001100011011110011000;
filter5[3][833] = 35'b11111110110011010010100101100100000;
filter5[3][834] = 35'b11111111011101100101010000111010000;
filter5[3][835] = 35'b00000000010000100101001101111011100;
filter5[3][836] = 35'b11111111010110010100111110000111000;
filter5[3][837] = 35'b11111101110111000111000000101100000;
filter5[3][838] = 35'b11111110011110110010011110110010000;
filter5[3][839] = 35'b11111110011101100101101100101010000;
filter5[3][840] = 35'b11111110010000111111010100100010000;
filter5[3][841] = 35'b11111101110111111000100110011100000;
filter5[3][842] = 35'b00000010000010101010010110011100000;
filter5[3][843] = 35'b00000011000110011111101111011000000;
filter5[3][844] = 35'b11111111000001101101111010001101000;
filter5[3][845] = 35'b11111111100101110000100101100011100;
filter5[3][846] = 35'b11111110111110101010001011011010000;
filter5[3][847] = 35'b11111110011100110011000110010100000;
filter5[3][848] = 35'b11111100111101110011100011110100000;
filter5[3][849] = 35'b11111100110000100001010001001000000;
filter5[3][850] = 35'b00000000100011010010011011011010000;
filter5[3][851] = 35'b00000000110011110010101011100011000;
filter5[3][852] = 35'b11111110110101101001001000101110000;
filter5[3][853] = 35'b00000001101001010110101000110000000;
filter5[3][854] = 35'b11111111101000011011100101000100100;
filter5[3][855] = 35'b11111110001000110111101101101100000;
filter5[3][856] = 35'b11111110110100100000010001011110000;
filter5[3][857] = 35'b11111100100100011110001000010100000;
filter5[3][858] = 35'b00000011010101111110010001010000000;
filter5[3][859] = 35'b00000001110111101111001011101010000;
filter5[3][860] = 35'b11111101111111101000000111001000000;
filter5[3][861] = 35'b00000010110111000001011101011100000;
filter5[3][862] = 35'b11111111110011011111111001101100110;
filter5[3][863] = 35'b11111111011100000101100100111011000;
filter5[3][864] = 35'b11111111111000001100111011011101100;
filter5[3][865] = 35'b11111110010101001010010000011000000;
filter5[3][866] = 35'b11111110111111100010010011110100000;
filter5[3][867] = 35'b00000100101010010110010100001000000;
filter5[3][868] = 35'b11111111011010100101001110000110000;
filter5[3][869] = 35'b11111100100110000101011100001000000;
filter5[3][870] = 35'b11111111000111010001000000100100000;
filter5[3][871] = 35'b11111101100111000010100000000000000;
filter5[3][872] = 35'b00000000001000101111011110100110110;
filter5[3][873] = 35'b00000100000011111110111001010000000;
filter5[3][874] = 35'b11111111100100101110011001100101100;
filter5[3][875] = 35'b00000001110010101000011100011100000;
filter5[3][876] = 35'b11111111000010000101000000000000000;
filter5[3][877] = 35'b11111100110010010100100101110000000;
filter5[3][878] = 35'b11111101011000111010100001010000000;
filter5[3][879] = 35'b11111101100110010000100101101100000;
filter5[3][880] = 35'b11111111101010110010110100001011000;
filter5[3][881] = 35'b00000100000010010011111111010000000;
filter5[3][882] = 35'b00000000000010010101101101010111000;
filter5[3][883] = 35'b00000100100111111101111100101000000;
filter5[3][884] = 35'b11111101010100000000100111000000000;
filter5[3][885] = 35'b11111111111100001111101010101101011;
filter5[3][886] = 35'b11111001010010110000100100010000000;
filter5[3][887] = 35'b11111111011110101000011111001010000;
filter5[3][888] = 35'b11111111110000011011011010000001000;
filter5[3][889] = 35'b00000001110010011011000011011100000;
filter5[3][890] = 35'b11111110000010010111011101010100000;
filter5[3][891] = 35'b00000001010010010111100010111110000;
filter5[3][892] = 35'b11111111001110010011101010100001000;
filter5[3][893] = 35'b11111100010101000100000010100100000;
filter5[3][894] = 35'b11111100111101001001111010110000000;
filter5[3][895] = 35'b11111110011011001010111001111100000;
filter5[3][896] = 35'b11111010100101110011100001101000000;
filter5[3][897] = 35'b11111100001110000011000100000100000;
filter5[3][898] = 35'b00000101100101011000010010010000000;
filter5[3][899] = 35'b00000101111110000111010010011000000;
filter5[3][900] = 35'b00001000001010101011010101110000000;
filter5[3][901] = 35'b11111010101010101010010110101000000;
filter5[3][902] = 35'b11111011101000011101001101000000000;
filter5[3][903] = 35'b11111111000111000010100110110101000;
filter5[3][904] = 35'b11111101100110000110011001110000000;
filter5[3][905] = 35'b11111011100010111101101111001000000;
filter5[3][906] = 35'b00000001010001111100000001000010000;
filter5[3][907] = 35'b11111011111111000011010101010000000;
filter5[3][908] = 35'b00000011010010011011101000110000000;
filter5[3][909] = 35'b11110111010000101101111001100000000;
filter5[3][910] = 35'b00000001000100111011101000111010000;
filter5[3][911] = 35'b11111010101011101010111001010000000;
filter5[3][912] = 35'b00000000011100000010110001101001000;
filter5[3][913] = 35'b11111101101100001000110001001000000;
filter5[3][914] = 35'b00000000110100000110110101100110000;
filter5[3][915] = 35'b11111101001101001100110101110100000;
filter5[3][916] = 35'b00000000101111000110100110001110000;
filter5[3][917] = 35'b11111110100110110001101101100010000;
filter5[3][918] = 35'b11111000111100010101010001101000000;
filter5[3][919] = 35'b11110011100000000101001001000000000;
filter5[3][920] = 35'b00000000010111111100011011000000000;
filter5[3][921] = 35'b11111110110101011111101110011100000;
filter5[3][922] = 35'b00000001111011110111101110111010000;
filter5[3][923] = 35'b00000001100100000111001011001100000;
filter5[3][924] = 35'b00000000011010000111110101001101000;
filter5[3][925] = 35'b00000000011100101101001011010100000;
filter5[3][926] = 35'b00000000011011111110010000111000000;
filter5[3][927] = 35'b11111010010100011111011011001000000;
filter5[3][928] = 35'b00000101111110010011000110111000000;
filter5[3][929] = 35'b11111111001100010000001111010101000;
filter5[3][930] = 35'b11111100101010100111010110101100000;
filter5[3][931] = 35'b00000010101000000001010100100000000;
filter5[3][932] = 35'b11111110010101110110110010110110000;
filter5[3][933] = 35'b11111101110010001011101111110000000;
filter5[3][934] = 35'b00000001100101000010000000011010000;
filter5[3][935] = 35'b11111101100010001001011110110100000;
filter5[3][936] = 35'b11111101001110000111100110101100000;
filter5[3][937] = 35'b00000100100011101000010110101000000;
filter5[3][938] = 35'b11111110110011100000101110101000000;
filter5[3][939] = 35'b00000001100110001110011000101000000;
filter5[3][940] = 35'b11111111111110101011111110100101011;
filter5[3][941] = 35'b11111110110010100110011100111100000;
filter5[3][942] = 35'b00000000000111010101110011010010001;
filter5[3][943] = 35'b00000001010001000100000011111010000;
filter5[3][944] = 35'b11111111101011011101100111010011000;
filter5[3][945] = 35'b00000001110111011011010110101000000;
filter5[3][946] = 35'b00000001010000101010010110110010000;
filter5[3][947] = 35'b00000001111000010101011000110100000;
filter5[3][948] = 35'b11111111011101001011111110111110000;
filter5[3][949] = 35'b11111111001010101001100010110011000;
filter5[3][950] = 35'b11111111111010000001100000011111101;
filter5[3][951] = 35'b11111100001111111000001100100000000;
filter5[3][952] = 35'b11111101010111101111001110000100000;
filter5[3][953] = 35'b00000111011111000000100010011000000;
filter5[3][954] = 35'b11111101101001101001001101000100000;
filter5[3][955] = 35'b00000000110110100111111010000010000;
filter5[3][956] = 35'b11111111110101010100100101101111000;
filter5[3][957] = 35'b11111101000110011110011110111100000;
filter5[3][958] = 35'b00000000101101010110010011111011000;
filter5[3][959] = 35'b11101001101110000111001100100000000;
filter5[3][960] = 35'b11111111101101111101001110101110100;
filter5[3][961] = 35'b00000000100011001101010111100110000;
filter5[3][962] = 35'b00000011000000100110101010100000000;
filter5[3][963] = 35'b00000100101010000100110100100000000;
filter5[3][964] = 35'b00001000001011001001111011100000000;
filter5[3][965] = 35'b00000101111000001111110001010000000;
filter5[3][966] = 35'b11111000010011001000111011000000000;
filter5[3][967] = 35'b11111001111101100000100111100000000;
filter5[3][968] = 35'b11111001001111010010111100000000000;
filter5[3][969] = 35'b00000001001100110000100001011100000;
filter5[3][970] = 35'b00000001010100011011110100011000000;
filter5[3][971] = 35'b11111101111011011011111101111000000;
filter5[3][972] = 35'b11111110101000110011010101000100000;
filter5[3][973] = 35'b11111110100111100110100110101100000;
filter5[3][974] = 35'b00000001011101010101001000110000000;
filter5[3][975] = 35'b00000101000110011110100101000000000;
filter5[3][976] = 35'b00000000100011010010110010010111000;
filter5[3][977] = 35'b11111111110101110001001110001110000;
filter5[3][978] = 35'b00000001110010010000111100000100000;
filter5[3][979] = 35'b11111101011010010110111110011000000;
filter5[3][980] = 35'b11111111111010000100100011101110110;
filter5[3][981] = 35'b00000000101110101010010101101000000;
filter5[3][982] = 35'b11111111101111000111011101110000100;
filter5[3][983] = 35'b00000000101011100111111101011000000;
filter5[3][984] = 35'b00000000010101001000100111000100000;
filter5[3][985] = 35'b11111110111001111000010100011000000;
filter5[3][986] = 35'b00000000111010011011011000000010000;
filter5[3][987] = 35'b00000001101001111101100100101110000;
filter5[3][988] = 35'b00000011010111000110111010000100000;
filter5[3][989] = 35'b00000011101100001001101010101100000;
filter5[3][990] = 35'b00000010000101000001000101010100000;
filter5[3][991] = 35'b00000000100110111111010010010001000;
filter5[3][992] = 35'b11110111001110101111100110010000000;
filter5[3][993] = 35'b11111111010110111111111011010110000;
filter5[3][994] = 35'b00000010111001101110000001010100000;
filter5[3][995] = 35'b00000011110011000010010110001000000;
filter5[3][996] = 35'b00000000110101100111100000111110000;
filter5[3][997] = 35'b11111010100101011111110011001000000;
filter5[3][998] = 35'b11111011011101111101011111100000000;
filter5[3][999] = 35'b11111011010000000110111110111000000;
filter5[3][1000] = 35'b00000001101111001110000100101110000;
filter5[3][1001] = 35'b11111101001100100110100010001000000;
filter5[3][1002] = 35'b00000001010000010010001010101000000;
filter5[3][1003] = 35'b00000010100110000101001010110100000;
filter5[3][1004] = 35'b00000000000100110011000011101110101;
filter5[3][1005] = 35'b11111011111100011111010011110000000;
filter5[3][1006] = 35'b11110100001001111100101011110000000;
filter5[3][1007] = 35'b11110111001001100000100100100000000;
filter5[3][1008] = 35'b11110010000001110011001100110000000;
filter5[3][1009] = 35'b11111111100000011101011011101000000;
filter5[3][1010] = 35'b11111111111001011100000111101101101;
filter5[3][1011] = 35'b00000000000111110000100111001011110;
filter5[3][1012] = 35'b11111100001101101000000011101100000;
filter5[3][1013] = 35'b11111101110101000011100000010100000;
filter5[3][1014] = 35'b11111100101110101100011110010100000;
filter5[3][1015] = 35'b11111000010100001110000101101000000;
filter5[3][1016] = 35'b11110110110000000110011000110000000;
filter5[3][1017] = 35'b00000001111111100000101110000110000;
filter5[3][1018] = 35'b00000111010101011101101101011000000;
filter5[3][1019] = 35'b00000100100100110100110101101000000;
filter5[3][1020] = 35'b11111001001101101010011111001000000;
filter5[3][1021] = 35'b11111111010001000011011000010100000;
filter5[3][1022] = 35'b00000000000010110111101101001101110;
filter5[3][1023] = 35'b11111000110101110001100100010000000;
filter5[4][0] = 35'b11111101011011101010001100011100000;
filter5[4][1] = 35'b00000010100000001011000111000100000;
filter5[4][2] = 35'b11111111000001110111110111101000000;
filter5[4][3] = 35'b11111111101010001101110101000011000;
filter5[4][4] = 35'b11110101100001111000100100100000000;
filter5[4][5] = 35'b11111101011010100000010101101000000;
filter5[4][6] = 35'b00000000100011011000100011011101000;
filter5[4][7] = 35'b11111110001101110010100001000110000;
filter5[4][8] = 35'b00000100011000010111101000011000000;
filter5[4][9] = 35'b00000001000111011101111101011000000;
filter5[4][10] = 35'b00000000110000000011101111111111000;
filter5[4][11] = 35'b00000001110011110011111010010100000;
filter5[4][12] = 35'b00000000111101111111010000011000000;
filter5[4][13] = 35'b11111011100001011100111111100000000;
filter5[4][14] = 35'b11110110001010111011101110100000000;
filter5[4][15] = 35'b11110101101001101000111001110000000;
filter5[4][16] = 35'b11111011100101000011011010001000000;
filter5[4][17] = 35'b11111011000111110111000110111000000;
filter5[4][18] = 35'b00000000101101011111010110101111000;
filter5[4][19] = 35'b11111110111001001010100010101000000;
filter5[4][20] = 35'b00000011110000100001000011001100000;
filter5[4][21] = 35'b00000011010111100101010101001100000;
filter5[4][22] = 35'b11111000110000000110110100110000000;
filter5[4][23] = 35'b11111011010010010011100111110000000;
filter5[4][24] = 35'b11111110001110101100010011001000000;
filter5[4][25] = 35'b00000000111110011000001100010101000;
filter5[4][26] = 35'b00000010010100001111100000110100000;
filter5[4][27] = 35'b00000001100011110000100101100010000;
filter5[4][28] = 35'b00000010000110101100000100100000000;
filter5[4][29] = 35'b11111000101111000000010011001000000;
filter5[4][30] = 35'b11111100110000110001010110010000000;
filter5[4][31] = 35'b11111111111101101010101010110111111;
filter5[4][32] = 35'b00000000010100100000010111010011100;
filter5[4][33] = 35'b00000001110100111100101011111010000;
filter5[4][34] = 35'b00000000100110000010100111000111000;
filter5[4][35] = 35'b11111111010110011000111111100000000;
filter5[4][36] = 35'b11111010100000100100110011100000000;
filter5[4][37] = 35'b00000101011110011000010001011000000;
filter5[4][38] = 35'b00000010011101111010110111010000000;
filter5[4][39] = 35'b11111110100100100111100110000110000;
filter5[4][40] = 35'b00000000000101010111110101000001001;
filter5[4][41] = 35'b00000100011110101000100101011000000;
filter5[4][42] = 35'b11111100001111000011111110101000000;
filter5[4][43] = 35'b00000000001001111000111000110100010;
filter5[4][44] = 35'b11111110110001110101101110110000000;
filter5[4][45] = 35'b00000000001011001101111001101011000;
filter5[4][46] = 35'b00000100101111101010100000110000000;
filter5[4][47] = 35'b11111100110111100110100000010100000;
filter5[4][48] = 35'b00000101100011010000100110100000000;
filter5[4][49] = 35'b00000010010100001111000110001100000;
filter5[4][50] = 35'b11111010010100100010100111011000000;
filter5[4][51] = 35'b00000001000001000110001011000110000;
filter5[4][52] = 35'b11111000000110010011111100010000000;
filter5[4][53] = 35'b00000000000110010111000100111101100;
filter5[4][54] = 35'b11111000101100110101011010111000000;
filter5[4][55] = 35'b00000100111101000010010011000000000;
filter5[4][56] = 35'b11111111111000101010000110100010110;
filter5[4][57] = 35'b00000001101110011000110101111110000;
filter5[4][58] = 35'b11110111100000011111100011100000000;
filter5[4][59] = 35'b00000001000001010001100110100000000;
filter5[4][60] = 35'b11111011011010101100001001111000000;
filter5[4][61] = 35'b00000011001011100001010000011000000;
filter5[4][62] = 35'b00000111011011001110110110101000000;
filter5[4][63] = 35'b00000001001111011000110110110110000;
filter5[4][64] = 35'b00000000010100100101000000111000100;
filter5[4][65] = 35'b11111101101001000010110100110100000;
filter5[4][66] = 35'b11111111111110001111101010100111000;
filter5[4][67] = 35'b00000100010010000111111101101000000;
filter5[4][68] = 35'b00000001101000110100000011110110000;
filter5[4][69] = 35'b11111110011110000000110100011000000;
filter5[4][70] = 35'b11111100111011010001000000011000000;
filter5[4][71] = 35'b11111011110100001111110111010000000;
filter5[4][72] = 35'b00000000000110111100011000001011101;
filter5[4][73] = 35'b00000011001011000010100111100100000;
filter5[4][74] = 35'b00000010100010010100111111101000000;
filter5[4][75] = 35'b00000011110111011001001111100100000;
filter5[4][76] = 35'b00000010011100010011100100100100000;
filter5[4][77] = 35'b00000000010010111101110001010101100;
filter5[4][78] = 35'b11111110110010011101100100101000000;
filter5[4][79] = 35'b11111100001000010011001010011100000;
filter5[4][80] = 35'b00000011111011011000010100000100000;
filter5[4][81] = 35'b11111010111001010000110011010000000;
filter5[4][82] = 35'b00000001011000110011011011101100000;
filter5[4][83] = 35'b00000001111100100010111000011100000;
filter5[4][84] = 35'b00000000110011101010101011010001000;
filter5[4][85] = 35'b00000000111000100100100001000010000;
filter5[4][86] = 35'b11111111110101100000100110101001010;
filter5[4][87] = 35'b00000010011011000101110000000000000;
filter5[4][88] = 35'b11111111010110110011011000101111000;
filter5[4][89] = 35'b11111111110110111010110110011001000;
filter5[4][90] = 35'b00000100000010110001101101010000000;
filter5[4][91] = 35'b11111111110011011010111100001010100;
filter5[4][92] = 35'b11111101111110010000010110000000000;
filter5[4][93] = 35'b11111111110101000110101000111011000;
filter5[4][94] = 35'b11111111111000100011101011001001000;
filter5[4][95] = 35'b11111110100110110101010110001100000;
filter5[4][96] = 35'b00000011100010110110110001011100000;
filter5[4][97] = 35'b11111111001011000111000111110111000;
filter5[4][98] = 35'b00000001001000111001100101111110000;
filter5[4][99] = 35'b11111110100110010110111001110010000;
filter5[4][100] = 35'b11111101100111110111111101111100000;
filter5[4][101] = 35'b11111111000011011100000000100000000;
filter5[4][102] = 35'b11111111000111101011111110000100000;
filter5[4][103] = 35'b11111011110110111010100010010000000;
filter5[4][104] = 35'b00000001011000110100010000011100000;
filter5[4][105] = 35'b00000000010100001111111000011010000;
filter5[4][106] = 35'b11111110111100000000001101011010000;
filter5[4][107] = 35'b00000000011000011101000001010110000;
filter5[4][108] = 35'b11111101001000100001011010010100000;
filter5[4][109] = 35'b11111001011110100111011010001000000;
filter5[4][110] = 35'b11111110011100011101011111100110000;
filter5[4][111] = 35'b11111010001111011000010111101000000;
filter5[4][112] = 35'b00000011100101100100101110100100000;
filter5[4][113] = 35'b00000100110000111101011011111000000;
filter5[4][114] = 35'b11111111111001100101100000111110010;
filter5[4][115] = 35'b00000000111111110111111101110111000;
filter5[4][116] = 35'b11111111100011000101011010000001000;
filter5[4][117] = 35'b00000000011000110111110101100100100;
filter5[4][118] = 35'b11111110100100110101110011011010000;
filter5[4][119] = 35'b11111010010001001101010000100000000;
filter5[4][120] = 35'b00000001001001000000110110110110000;
filter5[4][121] = 35'b00000110000101010111110001001000000;
filter5[4][122] = 35'b00000010011101100111111010010000000;
filter5[4][123] = 35'b00000001101111001111111111100010000;
filter5[4][124] = 35'b11111101101011111000110110000000000;
filter5[4][125] = 35'b00000000010110101101111100110011000;
filter5[4][126] = 35'b11111010000111111001011011010000000;
filter5[4][127] = 35'b11111110100011011111011011010000000;
filter5[4][128] = 35'b11111110000110001001000101010100000;
filter5[4][129] = 35'b11111101010111010101010000000100000;
filter5[4][130] = 35'b00000111111111001111001010100000000;
filter5[4][131] = 35'b00001000101111101100000100000000000;
filter5[4][132] = 35'b00000110101110001011010011100000000;
filter5[4][133] = 35'b11110101000001011110110110110000000;
filter5[4][134] = 35'b11110001010101110101110000000000000;
filter5[4][135] = 35'b11101110000011000101001010000000000;
filter5[4][136] = 35'b00001011000000111011111010000000000;
filter5[4][137] = 35'b00000110001001100010100100110000000;
filter5[4][138] = 35'b11111111010010001000100001000101000;
filter5[4][139] = 35'b00000001011000010000000011011000000;
filter5[4][140] = 35'b00000000011001110111000100100111100;
filter5[4][141] = 35'b00000011000011010101010111101100000;
filter5[4][142] = 35'b00000001001000010010101001101000000;
filter5[4][143] = 35'b11111000010111011001110111100000000;
filter5[4][144] = 35'b11111101001110000101001001011000000;
filter5[4][145] = 35'b11111111100000010111110110010001000;
filter5[4][146] = 35'b00000011000111000010001100101000000;
filter5[4][147] = 35'b00000001101000011100001110000000000;
filter5[4][148] = 35'b11111111111000010010111011110011011;
filter5[4][149] = 35'b11111111110001101010010010111101100;
filter5[4][150] = 35'b00000000101001101011100100100100000;
filter5[4][151] = 35'b11110111101001010111010000000000000;
filter5[4][152] = 35'b00000000100110001101000001010011000;
filter5[4][153] = 35'b11111111001101001011000010000111000;
filter5[4][154] = 35'b00000001001111111001010001001010000;
filter5[4][155] = 35'b00000001111111000111011000011100000;
filter5[4][156] = 35'b00000000100100010001110001011110000;
filter5[4][157] = 35'b00000010001010010110101101110000000;
filter5[4][158] = 35'b11111110010100100101000010011010000;
filter5[4][159] = 35'b00000000010110101100101100111110100;
filter5[4][160] = 35'b11111111111001000111100101100110010;
filter5[4][161] = 35'b11111110000000100101111001010000000;
filter5[4][162] = 35'b11111111100011100001011011001000100;
filter5[4][163] = 35'b11111100111110100010110111000100000;
filter5[4][164] = 35'b11110100010101000101111000010000000;
filter5[4][165] = 35'b11111010010001011011100001100000000;
filter5[4][166] = 35'b11110110110101000000011011010000000;
filter5[4][167] = 35'b11110011100101110110010011110000000;
filter5[4][168] = 35'b11111101100001101001001001000000000;
filter5[4][169] = 35'b00000010101110000001101000110100000;
filter5[4][170] = 35'b00000011101111100001011101111000000;
filter5[4][171] = 35'b11111001001111000110110101110000000;
filter5[4][172] = 35'b11110100110111111100101000000000000;
filter5[4][173] = 35'b11110011100011010010111000100000000;
filter5[4][174] = 35'b11101100110010001101101100000000000;
filter5[4][175] = 35'b11110001100010001010110011110000000;
filter5[4][176] = 35'b00000110011100110101010110000000000;
filter5[4][177] = 35'b00000011100110110101100100110000000;
filter5[4][178] = 35'b11111101111101010100111111110000000;
filter5[4][179] = 35'b11111110101110010111110001111110000;
filter5[4][180] = 35'b11110001010000010010011010010000000;
filter5[4][181] = 35'b11101111101011101110110011000000000;
filter5[4][182] = 35'b11111001100000000101100011001000000;
filter5[4][183] = 35'b11101111001110000000111011100000000;
filter5[4][184] = 35'b11111100111001111001100000011000000;
filter5[4][185] = 35'b11111000100101000110000011111000000;
filter5[4][186] = 35'b11111111110001010101110010000001110;
filter5[4][187] = 35'b00000100001100011011000000101000000;
filter5[4][188] = 35'b11110011000100101111111110000000000;
filter5[4][189] = 35'b11110010000111110001111010110000000;
filter5[4][190] = 35'b11110100001111001011100111100000000;
filter5[4][191] = 35'b11111110110011010010001001001110000;
filter5[4][192] = 35'b00000011110111011000111010010100000;
filter5[4][193] = 35'b11111001100110110011010110111000000;
filter5[4][194] = 35'b00000001100011000011101011011110000;
filter5[4][195] = 35'b00000101001000011011010010110000000;
filter5[4][196] = 35'b11111111011101011100110010111010000;
filter5[4][197] = 35'b11110101001101111110010111010000000;
filter5[4][198] = 35'b11110111100000000011011011010000000;
filter5[4][199] = 35'b11101111010001101111000001000000000;
filter5[4][200] = 35'b00000000001100011001100000001010010;
filter5[4][201] = 35'b00001100001011111100101011110000000;
filter5[4][202] = 35'b00000101001111111010000010100000000;
filter5[4][203] = 35'b00000100110111100101101010111000000;
filter5[4][204] = 35'b00001101010000101000001110000000000;
filter5[4][205] = 35'b00000101000011001110001010111000000;
filter5[4][206] = 35'b11111100000100110111010010111000000;
filter5[4][207] = 35'b11111000011100001001101100010000000;
filter5[4][208] = 35'b00001000001111011111010010110000000;
filter5[4][209] = 35'b00000001011000011111000110000110000;
filter5[4][210] = 35'b11111111111100101100011010011110010;
filter5[4][211] = 35'b00000010001000111011101111110100000;
filter5[4][212] = 35'b00000001000101110010001011100010000;
filter5[4][213] = 35'b00000000010111000101110010001110100;
filter5[4][214] = 35'b11111100001010101111000100101000000;
filter5[4][215] = 35'b11101101100001101011100001000000000;
filter5[4][216] = 35'b00001000110000001010000100100000000;
filter5[4][217] = 35'b11111101000110011110100111100000000;
filter5[4][218] = 35'b00000000001100001001111010110010010;
filter5[4][219] = 35'b00000011100111001000110000100100000;
filter5[4][220] = 35'b00000000011111000100100111111001000;
filter5[4][221] = 35'b11111100101100101010010101100000000;
filter5[4][222] = 35'b11111110001101001000000010011110000;
filter5[4][223] = 35'b11111111010110000101110100101010000;
filter5[4][224] = 35'b00001010000010011000011001110000000;
filter5[4][225] = 35'b00000101110111110000101000101000000;
filter5[4][226] = 35'b11111101111111100000100100100100000;
filter5[4][227] = 35'b00000001010101001010111100110000000;
filter5[4][228] = 35'b11111110110011011110101111101000000;
filter5[4][229] = 35'b11111111010000001100100001111010000;
filter5[4][230] = 35'b00000000101100010100001001101010000;
filter5[4][231] = 35'b11111100000110101000000011010100000;
filter5[4][232] = 35'b00000100000111100000001000111000000;
filter5[4][233] = 35'b00000000111000110001001100100010000;
filter5[4][234] = 35'b11111110110000101111100110100000000;
filter5[4][235] = 35'b11111111111111101000010010111100011;
filter5[4][236] = 35'b00000011111010110111000100011100000;
filter5[4][237] = 35'b11111111001000100110101110010110000;
filter5[4][238] = 35'b11111110101011110000101111100010000;
filter5[4][239] = 35'b11111111101000001011100010001110100;
filter5[4][240] = 35'b00000010001000011010111010010100000;
filter5[4][241] = 35'b11111101010010110110011010101000000;
filter5[4][242] = 35'b00000010110000001011011111110000000;
filter5[4][243] = 35'b00000000110111101000011110100000000;
filter5[4][244] = 35'b11111111111100001001010001111111011;
filter5[4][245] = 35'b11111111000010110000000000101110000;
filter5[4][246] = 35'b11111111111010000011011000000001010;
filter5[4][247] = 35'b11111111100001111101111111010111000;
filter5[4][248] = 35'b11111100111001101101010001101000000;
filter5[4][249] = 35'b00000010011001110011100010100100000;
filter5[4][250] = 35'b00000100010100111011011000011000000;
filter5[4][251] = 35'b11111111110100011011001100000110110;
filter5[4][252] = 35'b11111110111111011111001011110010000;
filter5[4][253] = 35'b11111110001000110101100100011100000;
filter5[4][254] = 35'b11111111000110110111110011011001000;
filter5[4][255] = 35'b11111110100110101111001011001110000;
filter5[4][256] = 35'b11111100111100001011101111000000000;
filter5[4][257] = 35'b11111100111100001100010000110100000;
filter5[4][258] = 35'b00000111111111100010110000000000000;
filter5[4][259] = 35'b00000010100111100101101011010000000;
filter5[4][260] = 35'b00000000000111100000000101001011110;
filter5[4][261] = 35'b11111011011000110110101101010000000;
filter5[4][262] = 35'b11111100101001111001100111010000000;
filter5[4][263] = 35'b11111110011110110100110110011110000;
filter5[4][264] = 35'b00000110101100100100000011010000000;
filter5[4][265] = 35'b00000111001000000110011101101000000;
filter5[4][266] = 35'b00000010101111000111001001100000000;
filter5[4][267] = 35'b00001001001001010101110100010000000;
filter5[4][268] = 35'b00001010000001000010001011010000000;
filter5[4][269] = 35'b11111110000001011001111111001000000;
filter5[4][270] = 35'b11111010001010101100000101111000000;
filter5[4][271] = 35'b11111011111010010011000110101000000;
filter5[4][272] = 35'b00000011110100010001101101010000000;
filter5[4][273] = 35'b00000010100111100100000000111100000;
filter5[4][274] = 35'b00000000101001110101000010100001000;
filter5[4][275] = 35'b00000000110110100111110100100100000;
filter5[4][276] = 35'b11111100111110000101001000110100000;
filter5[4][277] = 35'b11111111110111100011101101100001000;
filter5[4][278] = 35'b11111111100000001111110110101000000;
filter5[4][279] = 35'b11111001110000110111110100010000000;
filter5[4][280] = 35'b11111111101111010100110111000010000;
filter5[4][281] = 35'b11111101001101100110100000000000000;
filter5[4][282] = 35'b11111111110000110101001011000010010;
filter5[4][283] = 35'b00000011000010100110010001100100000;
filter5[4][284] = 35'b11111110111000110010011010000000000;
filter5[4][285] = 35'b00000000110111010110010011100001000;
filter5[4][286] = 35'b11111101100100100000001110111100000;
filter5[4][287] = 35'b11110110011011011101101111010000000;
filter5[4][288] = 35'b00000111110110011000111000010000000;
filter5[4][289] = 35'b00000000000111110010010100111111001;
filter5[4][290] = 35'b11111100010010101010001010000000000;
filter5[4][291] = 35'b00000011110110011001100101001000000;
filter5[4][292] = 35'b00000000001100011100010001100101110;
filter5[4][293] = 35'b11111101111101011011001000101100000;
filter5[4][294] = 35'b11111100010110111010111100111000000;
filter5[4][295] = 35'b11111001101011111100111100110000000;
filter5[4][296] = 35'b00000000101100011101011000011000000;
filter5[4][297] = 35'b00000010000010111010101011111100000;
filter5[4][298] = 35'b11111111001111011010011001001110000;
filter5[4][299] = 35'b00000010000101101110011111110100000;
filter5[4][300] = 35'b11111111001000110000011111100001000;
filter5[4][301] = 35'b11111111000000110001010011101100000;
filter5[4][302] = 35'b11111111011011010111001011101101000;
filter5[4][303] = 35'b11111110100000101001001000010000000;
filter5[4][304] = 35'b11111101001011100011101010011100000;
filter5[4][305] = 35'b00000001110001101101010111000010000;
filter5[4][306] = 35'b11111110001101111100011101110010000;
filter5[4][307] = 35'b11111111110100110001001111110011110;
filter5[4][308] = 35'b00000001011100000100110011110100000;
filter5[4][309] = 35'b00000000100010110010011001001001000;
filter5[4][310] = 35'b11111111111111000001110101110011100;
filter5[4][311] = 35'b11111011110101010100001010100000000;
filter5[4][312] = 35'b00001010110010111101100101110000000;
filter5[4][313] = 35'b00000101101110010111001110110000000;
filter5[4][314] = 35'b11111100111010111110010101001100000;
filter5[4][315] = 35'b00000010000011111011101101011000000;
filter5[4][316] = 35'b11111111001011100111101011100101000;
filter5[4][317] = 35'b00000001110101110101010000110010000;
filter5[4][318] = 35'b11111011110001111101011111101000000;
filter5[4][319] = 35'b11111000100011000111011100010000000;
filter5[4][320] = 35'b00000001111111100001011000010000000;
filter5[4][321] = 35'b11111110100100010000101100111000000;
filter5[4][322] = 35'b00000100110111101000110011111000000;
filter5[4][323] = 35'b00001001110101110101110000000000000;
filter5[4][324] = 35'b00000010000111011111000001000100000;
filter5[4][325] = 35'b11110110001101101011011101100000000;
filter5[4][326] = 35'b11111010101011111011101000110000000;
filter5[4][327] = 35'b11110011111110001000101100100000000;
filter5[4][328] = 35'b00000001100101010011111001111100000;
filter5[4][329] = 35'b00000010100101101110011010100000000;
filter5[4][330] = 35'b00000100100000010010011100010000000;
filter5[4][331] = 35'b00000001011110011101100001101000000;
filter5[4][332] = 35'b00000011101001011001000111101100000;
filter5[4][333] = 35'b11111111101010100000100010001010100;
filter5[4][334] = 35'b11111000001001000111000100000000000;
filter5[4][335] = 35'b11110011001110001010010111110000000;
filter5[4][336] = 35'b11111101100111100010010110000000000;
filter5[4][337] = 35'b11111110100011101101110110101110000;
filter5[4][338] = 35'b00000001010000001011011010111100000;
filter5[4][339] = 35'b11111111000101011110000001000111000;
filter5[4][340] = 35'b00000000110101110111011000101110000;
filter5[4][341] = 35'b00000001011001111111001011001010000;
filter5[4][342] = 35'b11111101000100011010011001000000000;
filter5[4][343] = 35'b11111101000011100101111111100100000;
filter5[4][344] = 35'b11111110011000011110010001011000000;
filter5[4][345] = 35'b00000011001000100010101101101000000;
filter5[4][346] = 35'b00000010110100101100011001111100000;
filter5[4][347] = 35'b11111100110101100001011101010100000;
filter5[4][348] = 35'b11111111011110010101011011100010000;
filter5[4][349] = 35'b11111011100001000011001011110000000;
filter5[4][350] = 35'b11111011111101101000111001111000000;
filter5[4][351] = 35'b00000100001101110110001110000000000;
filter5[4][352] = 35'b00000000001110000001111010110001000;
filter5[4][353] = 35'b00000111110001011000101100011000000;
filter5[4][354] = 35'b00000001000001001010110001010010000;
filter5[4][355] = 35'b11111111111011100110101111110011011;
filter5[4][356] = 35'b11111111011001101000111011011001000;
filter5[4][357] = 35'b11111101101010010111010010001100000;
filter5[4][358] = 35'b11111101010000110101110100000100000;
filter5[4][359] = 35'b11111111001001100001101110101010000;
filter5[4][360] = 35'b11111111010111101010000100000001000;
filter5[4][361] = 35'b00000100101010101000010000110000000;
filter5[4][362] = 35'b11111100000001111101101000111000000;
filter5[4][363] = 35'b11111101001110001101100101110100000;
filter5[4][364] = 35'b00000011100100111111011011101000000;
filter5[4][365] = 35'b11111111001000101000000101100000000;
filter5[4][366] = 35'b11111110010011111111101001111010000;
filter5[4][367] = 35'b00000000001010111011010011011001000;
filter5[4][368] = 35'b00000001111111000010001001001000000;
filter5[4][369] = 35'b00000010101001111011010101110100000;
filter5[4][370] = 35'b00000001001011011011111010001110000;
filter5[4][371] = 35'b11111110011011101011111001010110000;
filter5[4][372] = 35'b00000000001001010010101110011011110;
filter5[4][373] = 35'b00000000000101011110110001010110100;
filter5[4][374] = 35'b11111101101110111111001001001100000;
filter5[4][375] = 35'b00000010110000100010001011100100000;
filter5[4][376] = 35'b11111011111101000110001111011000000;
filter5[4][377] = 35'b00000001000100100101101001101100000;
filter5[4][378] = 35'b00000001100001010111011100111100000;
filter5[4][379] = 35'b11111110111001100110111111010000000;
filter5[4][380] = 35'b11111110100000011010111001011110000;
filter5[4][381] = 35'b00000000011100110001000001100010100;
filter5[4][382] = 35'b00000010000100000010111101001100000;
filter5[4][383] = 35'b00000010000110001100110011001000000;
filter5[4][384] = 35'b11111111100110110110101011110100100;
filter5[4][385] = 35'b00000000000010001010101010011001010;
filter5[4][386] = 35'b00000000111110001011001000110010000;
filter5[4][387] = 35'b00000010110110000111011111100000000;
filter5[4][388] = 35'b00000011110010011111101011101100000;
filter5[4][389] = 35'b00000000001110100100111010110010100;
filter5[4][390] = 35'b00000000110010110000111010100010000;
filter5[4][391] = 35'b00000010111010100001100010101000000;
filter5[4][392] = 35'b11111110001010101011101010011010000;
filter5[4][393] = 35'b00000010100110010010001101010000000;
filter5[4][394] = 35'b00000001100001110010001101001100000;
filter5[4][395] = 35'b00000101110110111101000111001000000;
filter5[4][396] = 35'b11111100000001001111110101000100000;
filter5[4][397] = 35'b11111101011100010101110111010100000;
filter5[4][398] = 35'b11111111000000010101000100111011000;
filter5[4][399] = 35'b11111111100111111111101110110101000;
filter5[4][400] = 35'b11111011000100101000001111000000000;
filter5[4][401] = 35'b11111101100010010010100111111000000;
filter5[4][402] = 35'b00000000000110101010001010010110100;
filter5[4][403] = 35'b00000010000101100110110000100000000;
filter5[4][404] = 35'b11111101100010011011111000100100000;
filter5[4][405] = 35'b11111110001001101011011001101000000;
filter5[4][406] = 35'b11111111111011001110011101010111100;
filter5[4][407] = 35'b11111110001010010110100111001110000;
filter5[4][408] = 35'b11111101000111110001010111000000000;
filter5[4][409] = 35'b11111100110111000011110110011100000;
filter5[4][410] = 35'b11111101010011101100011101011100000;
filter5[4][411] = 35'b11111101100010000001010011001100000;
filter5[4][412] = 35'b11111111011111010100001000010000000;
filter5[4][413] = 35'b00000000011100110000010110100110100;
filter5[4][414] = 35'b11111101001100000110010010001000000;
filter5[4][415] = 35'b11111011010100101000100100111000000;
filter5[4][416] = 35'b11111110101001100010000011010100000;
filter5[4][417] = 35'b00000000101111111111000101110101000;
filter5[4][418] = 35'b11111010111110111100011110000000000;
filter5[4][419] = 35'b00000000110111010011101000011101000;
filter5[4][420] = 35'b00000001010001111101001110101100000;
filter5[4][421] = 35'b11111011001010010000001110000000000;
filter5[4][422] = 35'b11111111110001101011101010101011010;
filter5[4][423] = 35'b11111110001001001011100011100010000;
filter5[4][424] = 35'b00000011010101101001110110100000000;
filter5[4][425] = 35'b11111011101111100011110101001000000;
filter5[4][426] = 35'b11111110111010000101110001101110000;
filter5[4][427] = 35'b11111001000101001011000011101000000;
filter5[4][428] = 35'b11111100110000101110011101100000000;
filter5[4][429] = 35'b00000001101100100110010100100010000;
filter5[4][430] = 35'b00000000110011000110010011101111000;
filter5[4][431] = 35'b00000001100110100100010110001100000;
filter5[4][432] = 35'b00000010110101111110011011010100000;
filter5[4][433] = 35'b00000001011111100111011111000110000;
filter5[4][434] = 35'b11111011011101000110101010111000000;
filter5[4][435] = 35'b11111111110111100011001011110010010;
filter5[4][436] = 35'b00000001000010010101010100110100000;
filter5[4][437] = 35'b00000011100101110010011010110100000;
filter5[4][438] = 35'b00000011011001000110100000100000000;
filter5[4][439] = 35'b00000010000100110001010110000100000;
filter5[4][440] = 35'b11111100110110001100001111101000000;
filter5[4][441] = 35'b11111010011011001110001101011000000;
filter5[4][442] = 35'b00000001101011000101101100001000000;
filter5[4][443] = 35'b00000001101011000001010010000110000;
filter5[4][444] = 35'b00000010001100100101111001010000000;
filter5[4][445] = 35'b00000010111111001010100101000000000;
filter5[4][446] = 35'b00001001110000111010110110110000000;
filter5[4][447] = 35'b00000011010110111110111001001100000;
filter5[4][448] = 35'b00000001100011011110110000001000000;
filter5[4][449] = 35'b00000000110010001100011000101110000;
filter5[4][450] = 35'b11111001110100101101000000011000000;
filter5[4][451] = 35'b11111000010100010010110000101000000;
filter5[4][452] = 35'b11111111100100001101100011100101000;
filter5[4][453] = 35'b11111111111000110000111010011111010;
filter5[4][454] = 35'b00000010010011110110110001101100000;
filter5[4][455] = 35'b11111110111101011110000010110010000;
filter5[4][456] = 35'b00000111000000000111101010101000000;
filter5[4][457] = 35'b00000001000010100111111101000110000;
filter5[4][458] = 35'b11111111011100011110001110011101000;
filter5[4][459] = 35'b00000100111010011001111110000000000;
filter5[4][460] = 35'b11111000001110100110101000001000000;
filter5[4][461] = 35'b11111100101001001110111100110100000;
filter5[4][462] = 35'b11111010000011111001111000000000000;
filter5[4][463] = 35'b00000010001111010110101011001100000;
filter5[4][464] = 35'b11111110110111100111110111010000000;
filter5[4][465] = 35'b11111010101101101100100100100000000;
filter5[4][466] = 35'b11111001110001010011101111000000000;
filter5[4][467] = 35'b11111010011111111001000110000000000;
filter5[4][468] = 35'b11110000101011101011000101000000000;
filter5[4][469] = 35'b11111100100010110001010011001000000;
filter5[4][470] = 35'b11111011111111101001110010011000000;
filter5[4][471] = 35'b11111010010000101011100111000000000;
filter5[4][472] = 35'b11101001011101001111000101000000000;
filter5[4][473] = 35'b11111000100111010111010101010000000;
filter5[4][474] = 35'b11111010101010010101001110110000000;
filter5[4][475] = 35'b11111110000110001000101000001110000;
filter5[4][476] = 35'b00000000001000111101000001101110000;
filter5[4][477] = 35'b11111110101011111000111000010110000;
filter5[4][478] = 35'b11111110001100110101011001001010000;
filter5[4][479] = 35'b00000010000000110001101001000100000;
filter5[4][480] = 35'b11111000101001110000110101110000000;
filter5[4][481] = 35'b11101101011011001100011001000000000;
filter5[4][482] = 35'b11111011000001111001010010100000000;
filter5[4][483] = 35'b11110111111111001011011001010000000;
filter5[4][484] = 35'b00000000011010000010110010111010100;
filter5[4][485] = 35'b00000011001111010110111001001000000;
filter5[4][486] = 35'b00000101011010011001010111100000000;
filter5[4][487] = 35'b00000001000110111000011000000000000;
filter5[4][488] = 35'b00000100000001011110001100011000000;
filter5[4][489] = 35'b00000000000001000011001000011010001;
filter5[4][490] = 35'b00000000000001100100001001000110101;
filter5[4][491] = 35'b11111011000010000110011101100000000;
filter5[4][492] = 35'b11111111011010000000111001111111000;
filter5[4][493] = 35'b11111011001011011001101010110000000;
filter5[4][494] = 35'b11111110101101110010100110100100000;
filter5[4][495] = 35'b11111101110011001010111000101100000;
filter5[4][496] = 35'b00000100010110111110000001101000000;
filter5[4][497] = 35'b00000010111111101000111000000100000;
filter5[4][498] = 35'b00000100110100110101101110011000000;
filter5[4][499] = 35'b11111110100110000110100111111000000;
filter5[4][500] = 35'b11111101011010100001110010001100000;
filter5[4][501] = 35'b11111001101001100110000010001000000;
filter5[4][502] = 35'b11111110101011100000011010100010000;
filter5[4][503] = 35'b00000000011100000011010001000011100;
filter5[4][504] = 35'b00000001111111100001100001000100000;
filter5[4][505] = 35'b11111111110101001110001011111000010;
filter5[4][506] = 35'b00000101001100011111010111100000000;
filter5[4][507] = 35'b00000001001010100110100101001000000;
filter5[4][508] = 35'b11111111101010110000011101100000100;
filter5[4][509] = 35'b11111100000111111000110100001100000;
filter5[4][510] = 35'b00000101101011000010000001110000000;
filter5[4][511] = 35'b00000010000001100111011101101000000;
filter5[4][512] = 35'b00000001000000111100011111000100000;
filter5[4][513] = 35'b00000100010100010100001100011000000;
filter5[4][514] = 35'b00000001011101001010000001010000000;
filter5[4][515] = 35'b11111111101110001100110100011101100;
filter5[4][516] = 35'b00000111101110101001110111011000000;
filter5[4][517] = 35'b11111100010100010111101111001100000;
filter5[4][518] = 35'b11111101000010100010001010111000000;
filter5[4][519] = 35'b00000010011011010110001001101000000;
filter5[4][520] = 35'b00000000010100111100001110110000100;
filter5[4][521] = 35'b00000001001100000101110110001000000;
filter5[4][522] = 35'b00000010001110011010011101101100000;
filter5[4][523] = 35'b00000010111100111101111000110100000;
filter5[4][524] = 35'b11111011111101010110000110101000000;
filter5[4][525] = 35'b00000001000110000111111011111100000;
filter5[4][526] = 35'b11111111101010111111100100100000000;
filter5[4][527] = 35'b11111011100001100001100100110000000;
filter5[4][528] = 35'b00000000001000100011110100001000000;
filter5[4][529] = 35'b11111111110010101110100111111110010;
filter5[4][530] = 35'b00000000010101110011001100110001000;
filter5[4][531] = 35'b11111110001000110111110011001100000;
filter5[4][532] = 35'b00000000111100100111010010010100000;
filter5[4][533] = 35'b00000000001110000101111010110011100;
filter5[4][534] = 35'b11111110011101111011001100111110000;
filter5[4][535] = 35'b11111111010011001110011101100101000;
filter5[4][536] = 35'b00000010111111010010001000110100000;
filter5[4][537] = 35'b00000000010110101111111100011110100;
filter5[4][538] = 35'b00000001001100011110110001111010000;
filter5[4][539] = 35'b11111110110100110111000000111100000;
filter5[4][540] = 35'b00000001100100001000110011100110000;
filter5[4][541] = 35'b00000001001011011111110000110010000;
filter5[4][542] = 35'b00000000000110011111110001000010111;
filter5[4][543] = 35'b11111101100011000000100111001100000;
filter5[4][544] = 35'b11111101111110010101001111010100000;
filter5[4][545] = 35'b00000001101101000010010000100100000;
filter5[4][546] = 35'b11111100101110101111111111011000000;
filter5[4][547] = 35'b00000001001110110101010100000010000;
filter5[4][548] = 35'b00000001011101011110011010110000000;
filter5[4][549] = 35'b00000000001100001011100000101111000;
filter5[4][550] = 35'b11111011101001010000111110101000000;
filter5[4][551] = 35'b00000000110110110110011100010001000;
filter5[4][552] = 35'b00000011111010001110000110001000000;
filter5[4][553] = 35'b11111110111010000100011001011000000;
filter5[4][554] = 35'b11111001101011011110101000110000000;
filter5[4][555] = 35'b00000001110011000101001011100100000;
filter5[4][556] = 35'b11111110000010010010001010000110000;
filter5[4][557] = 35'b11111111101111100010101101100010100;
filter5[4][558] = 35'b00000001100000001011010011011010000;
filter5[4][559] = 35'b11111110111000111100100110110100000;
filter5[4][560] = 35'b00000011001000011010101001011000000;
filter5[4][561] = 35'b11111010110101100110111101000000000;
filter5[4][562] = 35'b00000010111100100110101011111100000;
filter5[4][563] = 35'b00000001000110000111000001101010000;
filter5[4][564] = 35'b11111111101000010100010000111100000;
filter5[4][565] = 35'b11111111011011011100000011000111000;
filter5[4][566] = 35'b11111111100100010101000110010100000;
filter5[4][567] = 35'b11111011000111111010011001010000000;
filter5[4][568] = 35'b00000100010111001010011111010000000;
filter5[4][569] = 35'b11111010011000000110010100111000000;
filter5[4][570] = 35'b11111101111001100101110110101000000;
filter5[4][571] = 35'b11111111110000011111101000111100110;
filter5[4][572] = 35'b11111111011011110111000110110111000;
filter5[4][573] = 35'b00000010011001001010011000110000000;
filter5[4][574] = 35'b00000001110011000110000100111010000;
filter5[4][575] = 35'b00000000110001100100011011111101000;
filter5[4][576] = 35'b00000001000010101101000100011010000;
filter5[4][577] = 35'b00000001010011011111100111010100000;
filter5[4][578] = 35'b11111111001110100011101101111110000;
filter5[4][579] = 35'b11111110100110100110101011010100000;
filter5[4][580] = 35'b00001001001110110111111010000000000;
filter5[4][581] = 35'b11111101100100111100011110000000000;
filter5[4][582] = 35'b11111001111100001110111001010000000;
filter5[4][583] = 35'b00000000001110000011101011011101000;
filter5[4][584] = 35'b11110101101001101110001100000000000;
filter5[4][585] = 35'b00000000001111111111010000101110110;
filter5[4][586] = 35'b00000001001001110001010110100110000;
filter5[4][587] = 35'b00001000000010100111010011100000000;
filter5[4][588] = 35'b11111100001100110101100110100100000;
filter5[4][589] = 35'b00000001110001011000110010000000000;
filter5[4][590] = 35'b11111110101001011100001111011010000;
filter5[4][591] = 35'b11111000000110000010000010100000000;
filter5[4][592] = 35'b11110110011101100100010010110000000;
filter5[4][593] = 35'b00000010111000010100001101100000000;
filter5[4][594] = 35'b00000001101010110001111010011110000;
filter5[4][595] = 35'b00000000011000111011011111101110100;
filter5[4][596] = 35'b00000001010110010100101001000110000;
filter5[4][597] = 35'b11111111010000001001000001110100000;
filter5[4][598] = 35'b00000000000001010111111111010001110;
filter5[4][599] = 35'b11111010010011101111110101010000000;
filter5[4][600] = 35'b11111110100110110001001110111000000;
filter5[4][601] = 35'b00000011010101000100010110100100000;
filter5[4][602] = 35'b00000001101001001110011010001010000;
filter5[4][603] = 35'b11111110111111000101011100001110000;
filter5[4][604] = 35'b11111110011011001110100110001000000;
filter5[4][605] = 35'b11111111011000000000101100111000000;
filter5[4][606] = 35'b00000001000011100100101111111000000;
filter5[4][607] = 35'b11111011100100111110101001100000000;
filter5[4][608] = 35'b11110101001001000111101111110000000;
filter5[4][609] = 35'b00000011111001001001010100101000000;
filter5[4][610] = 35'b11111111001001110100001010111101000;
filter5[4][611] = 35'b00000000100001000010110101100111000;
filter5[4][612] = 35'b11111110001110011111000001111100000;
filter5[4][613] = 35'b11111110101001100101010110010010000;
filter5[4][614] = 35'b11111110110010000010011001110000000;
filter5[4][615] = 35'b11111110111100110111011101011100000;
filter5[4][616] = 35'b11111100000010101001011011000000000;
filter5[4][617] = 35'b11111100000001100011010011110100000;
filter5[4][618] = 35'b00000001001011000110111100011010000;
filter5[4][619] = 35'b00000000010000010011100111001000000;
filter5[4][620] = 35'b00000000011111011111000011000110000;
filter5[4][621] = 35'b11111110101011010110100110000000000;
filter5[4][622] = 35'b00000001000000001011100011011000000;
filter5[4][623] = 35'b00000000111111001111110000011001000;
filter5[4][624] = 35'b11111101111100001011111000001100000;
filter5[4][625] = 35'b11111101001010010000101110101000000;
filter5[4][626] = 35'b00000100000110110111000101011000000;
filter5[4][627] = 35'b00000001001011010011110011111010000;
filter5[4][628] = 35'b00000001111101110111111010111000000;
filter5[4][629] = 35'b11111101010110011001011011100000000;
filter5[4][630] = 35'b11111101100110001100000111111100000;
filter5[4][631] = 35'b00000001001100000011100000001100000;
filter5[4][632] = 35'b11111110010010011101100011100000000;
filter5[4][633] = 35'b11111110001000110001000101100110000;
filter5[4][634] = 35'b00000010001111111101010111100000000;
filter5[4][635] = 35'b00000001100101111110000101010010000;
filter5[4][636] = 35'b00000001101110011010100011001010000;
filter5[4][637] = 35'b11111111100111000010000110110110000;
filter5[4][638] = 35'b11111111001111000111101111000111000;
filter5[4][639] = 35'b00000000000000000110111101101110001;
filter5[4][640] = 35'b11111001001011101111110001100000000;
filter5[4][641] = 35'b00000001011000101001101100000000000;
filter5[4][642] = 35'b11111110101000110111111110110110000;
filter5[4][643] = 35'b11111110100001110101111110101010000;
filter5[4][644] = 35'b11111111100000001011010000100101000;
filter5[4][645] = 35'b11111001101110000000011000110000000;
filter5[4][646] = 35'b00000001101101011100100100100010000;
filter5[4][647] = 35'b00000000011100011000101101010111100;
filter5[4][648] = 35'b11111111111111100010001010010100101;
filter5[4][649] = 35'b00001001001101010000100100110000000;
filter5[4][650] = 35'b11111001101111100110001011101000000;
filter5[4][651] = 35'b11111101111100011111110001011100000;
filter5[4][652] = 35'b11111100011001000011111010001000000;
filter5[4][653] = 35'b00000011001001000111111001000100000;
filter5[4][654] = 35'b11111111000010110110000001101100000;
filter5[4][655] = 35'b11111011010000010101101010100000000;
filter5[4][656] = 35'b11110111101000111010101100100000000;
filter5[4][657] = 35'b11111010110100000011000001100000000;
filter5[4][658] = 35'b00000001100001101110101111010110000;
filter5[4][659] = 35'b00000011011101101001101000000000000;
filter5[4][660] = 35'b00000011001000100001101101001000000;
filter5[4][661] = 35'b11111011110011111010111011010000000;
filter5[4][662] = 35'b00000010111011001001110111111000000;
filter5[4][663] = 35'b11110101110100110101111100010000000;
filter5[4][664] = 35'b11110111111010011100000110100000000;
filter5[4][665] = 35'b11110111111111111111110011100000000;
filter5[4][666] = 35'b00000011011110001011011101000000000;
filter5[4][667] = 35'b00000011010111010001101111111100000;
filter5[4][668] = 35'b00000000101111011010111101011110000;
filter5[4][669] = 35'b11111111111101001101111001001100110;
filter5[4][670] = 35'b11111110010011010010110111010100000;
filter5[4][671] = 35'b11111010110010101101011110100000000;
filter5[4][672] = 35'b11111001011110001100110110010000000;
filter5[4][673] = 35'b00000001011100010110100111111000000;
filter5[4][674] = 35'b11110111111110101010110101100000000;
filter5[4][675] = 35'b00000000101000011100101011100001000;
filter5[4][676] = 35'b00000010001011011110001000100100000;
filter5[4][677] = 35'b00000000101010110011000101101100000;
filter5[4][678] = 35'b00000010001011010000010111010100000;
filter5[4][679] = 35'b00000011001011011110110000100100000;
filter5[4][680] = 35'b11111100110011001100100110111000000;
filter5[4][681] = 35'b11111001110011010011101011001000000;
filter5[4][682] = 35'b11111001101010111000101100000000000;
filter5[4][683] = 35'b11111111000101110010100011111111000;
filter5[4][684] = 35'b00000001000001000010111001010100000;
filter5[4][685] = 35'b00000000101111100000001100010100000;
filter5[4][686] = 35'b11111111001001010101110110110101000;
filter5[4][687] = 35'b11111110101000000101110000100000000;
filter5[4][688] = 35'b00000011100110110111101111001100000;
filter5[4][689] = 35'b00000010010000011001110110101000000;
filter5[4][690] = 35'b00000001110101000101010101101000000;
filter5[4][691] = 35'b11111110111011110101010101000110000;
filter5[4][692] = 35'b11111101111011010001111000000000000;
filter5[4][693] = 35'b11111010110111100101100001101000000;
filter5[4][694] = 35'b00000001110111111001001010011000000;
filter5[4][695] = 35'b11111111000111000000010101010011000;
filter5[4][696] = 35'b00000011000011010100011011100000000;
filter5[4][697] = 35'b11111110111100010100101011100000000;
filter5[4][698] = 35'b00000010001011101110111101010100000;
filter5[4][699] = 35'b11111111100000010100101101101010000;
filter5[4][700] = 35'b11111011110000000000001000101000000;
filter5[4][701] = 35'b00000100111001111111101001001000000;
filter5[4][702] = 35'b00000101100100011101010011010000000;
filter5[4][703] = 35'b00000000001001101000101010010000100;
filter5[4][704] = 35'b11111101101111111101001000000100000;
filter5[4][705] = 35'b11111101000010000110100010111100000;
filter5[4][706] = 35'b00000001001001110001111000011100000;
filter5[4][707] = 35'b00000000111100111100101001000111000;
filter5[4][708] = 35'b11111111101110101010110101010010000;
filter5[4][709] = 35'b11111100101110000100110000001100000;
filter5[4][710] = 35'b11111110100001011111110001111000000;
filter5[4][711] = 35'b11111110110000001100000110001100000;
filter5[4][712] = 35'b11111110001010111101101011111110000;
filter5[4][713] = 35'b11111100010100010101001101111100000;
filter5[4][714] = 35'b11111111110110111110111100000010000;
filter5[4][715] = 35'b11111110110011011001011000010100000;
filter5[4][716] = 35'b00000010111110011001100111011000000;
filter5[4][717] = 35'b11111111010110101101001011101111000;
filter5[4][718] = 35'b11111101100010011110001000001000000;
filter5[4][719] = 35'b11111111010010010001100001001110000;
filter5[4][720] = 35'b00000010000111001111001100100100000;
filter5[4][721] = 35'b11111101010011110001000001100100000;
filter5[4][722] = 35'b00000000010001110100111001011010100;
filter5[4][723] = 35'b00000010011110001111100001110100000;
filter5[4][724] = 35'b00000000111001110110010101001100000;
filter5[4][725] = 35'b00000001110100011011000111010100000;
filter5[4][726] = 35'b11111100011101100010011001100100000;
filter5[4][727] = 35'b11111011101011100100100101111000000;
filter5[4][728] = 35'b00000011001100010011000011000100000;
filter5[4][729] = 35'b11111110111110100110000011101010000;
filter5[4][730] = 35'b00000011000000100001001001100000000;
filter5[4][731] = 35'b00000001001000111110000001101010000;
filter5[4][732] = 35'b00000010011010011000110101011000000;
filter5[4][733] = 35'b11111101100110100101000101110000000;
filter5[4][734] = 35'b11111111111010101011110011111010011;
filter5[4][735] = 35'b11111101101000110000111010100100000;
filter5[4][736] = 35'b00000011110110011010110010111000000;
filter5[4][737] = 35'b00000000001010110000001000000101110;
filter5[4][738] = 35'b11111110010011100000101011111100000;
filter5[4][739] = 35'b00000001000010101100001000010110000;
filter5[4][740] = 35'b00000000001011110110011110000110010;
filter5[4][741] = 35'b11111110101100001100110101101110000;
filter5[4][742] = 35'b00000000011110100101011101011110000;
filter5[4][743] = 35'b11111011010010010100001011111000000;
filter5[4][744] = 35'b00000000111100101010001100011100000;
filter5[4][745] = 35'b00000011110111111111101010111000000;
filter5[4][746] = 35'b11111111011110001010101000110010000;
filter5[4][747] = 35'b11111111011100100000111000111011000;
filter5[4][748] = 35'b00000000101110010101100011011001000;
filter5[4][749] = 35'b11111100111101011000110110010100000;
filter5[4][750] = 35'b11111101111111010111011101100000000;
filter5[4][751] = 35'b11111110110101010010100011101000000;
filter5[4][752] = 35'b00000001011111010000011100001110000;
filter5[4][753] = 35'b00000000100100101111111011100110000;
filter5[4][754] = 35'b00000010001100001000001010011000000;
filter5[4][755] = 35'b00000001101111110001010000010100000;
filter5[4][756] = 35'b11111111110000001001101010100110000;
filter5[4][757] = 35'b11111110100010100101010101010000000;
filter5[4][758] = 35'b11111101011111010000000100100000000;
filter5[4][759] = 35'b11111110011101000000110000000000000;
filter5[4][760] = 35'b11111111011000001000110011111111000;
filter5[4][761] = 35'b00000000100001000111001011001001000;
filter5[4][762] = 35'b00000010111000101111100011010000000;
filter5[4][763] = 35'b00000001101110001101010011100000000;
filter5[4][764] = 35'b11111111101100100001110110100110000;
filter5[4][765] = 35'b11111110000001000111001111011000000;
filter5[4][766] = 35'b11111110111001100010000010111010000;
filter5[4][767] = 35'b11111101110101100011111110101100000;
filter5[4][768] = 35'b00000000001000011101010111001011010;
filter5[4][769] = 35'b00000010100010101001111110010100000;
filter5[4][770] = 35'b00000010111110010000100101100100000;
filter5[4][771] = 35'b00000010000111101011011101010000000;
filter5[4][772] = 35'b11111111011111000000010110101001000;
filter5[4][773] = 35'b11111111001011110001011110010000000;
filter5[4][774] = 35'b00000010000010011010000011001100000;
filter5[4][775] = 35'b00000010010011011010110011110100000;
filter5[4][776] = 35'b00000110111010110011100111101000000;
filter5[4][777] = 35'b00000010011010010111000011010000000;
filter5[4][778] = 35'b00000100111101011100011101001000000;
filter5[4][779] = 35'b11111001001000101100001101010000000;
filter5[4][780] = 35'b11111110111100101010010010001110000;
filter5[4][781] = 35'b11111111111110101100101011010011000;
filter5[4][782] = 35'b00000100111000010101101100011000000;
filter5[4][783] = 35'b11111111110010111001011011110000110;
filter5[4][784] = 35'b00000011100000110011001111101100000;
filter5[4][785] = 35'b00000011011110111010011101010100000;
filter5[4][786] = 35'b11111101010100110000100111100100000;
filter5[4][787] = 35'b11111101011011110001110010100100000;
filter5[4][788] = 35'b11110101110100101100111100100000000;
filter5[4][789] = 35'b11111001010011101101111111101000000;
filter5[4][790] = 35'b11111000101111100001001100010000000;
filter5[4][791] = 35'b00000101100001001001010110000000000;
filter5[4][792] = 35'b00000011101001010111001111110000000;
filter5[4][793] = 35'b00000100000111001010001000111000000;
filter5[4][794] = 35'b11111110001100100101100110100100000;
filter5[4][795] = 35'b11111001100111100011001110010000000;
filter5[4][796] = 35'b11111101000111011000001011000000000;
filter5[4][797] = 35'b11111010010010110100001110010000000;
filter5[4][798] = 35'b11111101011100100010111000000000000;
filter5[4][799] = 35'b00000001000001100110000100010110000;
filter5[4][800] = 35'b00000010010000011011000100001000000;
filter5[4][801] = 35'b11111011101011111101101011010000000;
filter5[4][802] = 35'b00000000000100001001000001000001111;
filter5[4][803] = 35'b11111000100011111110000111011000000;
filter5[4][804] = 35'b00000000100010100101100100101001000;
filter5[4][805] = 35'b11111111001010110000110010011110000;
filter5[4][806] = 35'b00000011001011110001001111000000000;
filter5[4][807] = 35'b11111011111000010001101110011000000;
filter5[4][808] = 35'b00000101110110001001000000010000000;
filter5[4][809] = 35'b11111111100110111110010110000100100;
filter5[4][810] = 35'b11110111100011110000000001110000000;
filter5[4][811] = 35'b11111010101011000001000111110000000;
filter5[4][812] = 35'b11111110110111100000110100101010000;
filter5[4][813] = 35'b00000010101001000011110011001000000;
filter5[4][814] = 35'b11111111101101001000001000000010000;
filter5[4][815] = 35'b00000000111110111111100111001011000;
filter5[4][816] = 35'b00000010100001110011001100001000000;
filter5[4][817] = 35'b11111110011001101100001010101010000;
filter5[4][818] = 35'b00000010000000100001100010110000000;
filter5[4][819] = 35'b11111111110101110001100111010000000;
filter5[4][820] = 35'b00000010111001101001001011011000000;
filter5[4][821] = 35'b11111110011110000100111011011000000;
filter5[4][822] = 35'b11111010101011111000111001100000000;
filter5[4][823] = 35'b00000011100111011000100000111000000;
filter5[4][824] = 35'b00000000110111110000100011000011000;
filter5[4][825] = 35'b11111100011110001010010101000000000;
filter5[4][826] = 35'b00000010100010101000000010101100000;
filter5[4][827] = 35'b00000001100100010000000011001110000;
filter5[4][828] = 35'b00000000010000001000101111011011000;
filter5[4][829] = 35'b11111110001111110011000111000010000;
filter5[4][830] = 35'b11111110001100000111011000110010000;
filter5[4][831] = 35'b00001000000011010110101000110000000;
filter5[4][832] = 35'b11111110100111101111101001010000000;
filter5[4][833] = 35'b11111101101111000000001100010100000;
filter5[4][834] = 35'b11111101010111001101011110101100000;
filter5[4][835] = 35'b11111111101100011101100010011110000;
filter5[4][836] = 35'b11111100111110101010001000101000000;
filter5[4][837] = 35'b11111110111011100011010011011010000;
filter5[4][838] = 35'b11111111000110100111101000011001000;
filter5[4][839] = 35'b11111111000100010101000011000110000;
filter5[4][840] = 35'b11111011111111000000111000110000000;
filter5[4][841] = 35'b11111111001110111110010101100100000;
filter5[4][842] = 35'b11111111111000111111101100101000100;
filter5[4][843] = 35'b00000001101111000011001101001110000;
filter5[4][844] = 35'b00000011100010000101001010010100000;
filter5[4][845] = 35'b11111111101110010011010011001100000;
filter5[4][846] = 35'b11111110100000010110100101101100000;
filter5[4][847] = 35'b11111110011010001110010000110010000;
filter5[4][848] = 35'b11111111100110110110011101000101000;
filter5[4][849] = 35'b00000001101001101100100000101110000;
filter5[4][850] = 35'b00000000011111000101101001001110100;
filter5[4][851] = 35'b00000001110100100001101001010000000;
filter5[4][852] = 35'b00000001010111011111001100111110000;
filter5[4][853] = 35'b11111111000010000000011010110011000;
filter5[4][854] = 35'b11111111001110000111110000101000000;
filter5[4][855] = 35'b11111100001100100111000100110000000;
filter5[4][856] = 35'b00000011110001000101100010011100000;
filter5[4][857] = 35'b11111111111011101011001100000001100;
filter5[4][858] = 35'b11111111000000101111001110110100000;
filter5[4][859] = 35'b00000001001101110100011000010100000;
filter5[4][860] = 35'b11111110100111100111111011000000000;
filter5[4][861] = 35'b00000001110101100010010111000100000;
filter5[4][862] = 35'b11111111011011111100001110000111000;
filter5[4][863] = 35'b11111111101010111110010100001110000;
filter5[4][864] = 35'b11111110101101100100101100111000000;
filter5[4][865] = 35'b11111111001100101100010111011011000;
filter5[4][866] = 35'b00000000011111011010111001011001000;
filter5[4][867] = 35'b11111111010110010101101101010111000;
filter5[4][868] = 35'b11111111010011111011011011011001000;
filter5[4][869] = 35'b00000001000010101111111000100110000;
filter5[4][870] = 35'b11111100010111101001110011010000000;
filter5[4][871] = 35'b11111011111110110100001011011000000;
filter5[4][872] = 35'b00000011010111111111110110110000000;
filter5[4][873] = 35'b11111111100111100101011010110000000;
filter5[4][874] = 35'b00000000101001011010110101100010000;
filter5[4][875] = 35'b00000011001111100011110001111100000;
filter5[4][876] = 35'b00000011111111011010111101100000000;
filter5[4][877] = 35'b11111110011110100010011001100000000;
filter5[4][878] = 35'b11111011111000011001010000010000000;
filter5[4][879] = 35'b11111000110100001010011000100000000;
filter5[4][880] = 35'b00000001001010010010010011100110000;
filter5[4][881] = 35'b00000010100001101100110010010100000;
filter5[4][882] = 35'b00000000100000101000011011101010000;
filter5[4][883] = 35'b11111110000110001101000100001000000;
filter5[4][884] = 35'b11111100001101000001111000101000000;
filter5[4][885] = 35'b11111010101110011100111111100000000;
filter5[4][886] = 35'b11111110101001100010010001011100000;
filter5[4][887] = 35'b11111011101010000001100000011000000;
filter5[4][888] = 35'b00000001110011011000011001110110000;
filter5[4][889] = 35'b00000101001000100100110111000000000;
filter5[4][890] = 35'b00000000101111000101001110010110000;
filter5[4][891] = 35'b00000010100001011011111100111000000;
filter5[4][892] = 35'b00000010001110111100110100110100000;
filter5[4][893] = 35'b11111100001010110100001001110000000;
filter5[4][894] = 35'b11111100100100101110111100001100000;
filter5[4][895] = 35'b11111100101010011000101011010000000;
filter5[4][896] = 35'b00000011001001001101011100101000000;
filter5[4][897] = 35'b00001001011001001110101100100000000;
filter5[4][898] = 35'b00001000011000110000001111100000000;
filter5[4][899] = 35'b00000110100100010101010000110000000;
filter5[4][900] = 35'b11111010000010011100110011100000000;
filter5[4][901] = 35'b11111011110110111110110100110000000;
filter5[4][902] = 35'b11111011100000111111101000111000000;
filter5[4][903] = 35'b11111000010011010100100010001000000;
filter5[4][904] = 35'b00000011101110000001111111100100000;
filter5[4][905] = 35'b00000010001010101001100101001000000;
filter5[4][906] = 35'b11111101101111011000111011001000000;
filter5[4][907] = 35'b11111111101010110101001111100010100;
filter5[4][908] = 35'b00000001111100011010010010111100000;
filter5[4][909] = 35'b00000000111000001000100110101000000;
filter5[4][910] = 35'b11111000011110001111101111110000000;
filter5[4][911] = 35'b11111011101101001010001011101000000;
filter5[4][912] = 35'b00000110010011100101001011100000000;
filter5[4][913] = 35'b11111110001011011001110100011100000;
filter5[4][914] = 35'b11111101101001000011111001011100000;
filter5[4][915] = 35'b00000000110110100101001100100011000;
filter5[4][916] = 35'b00000010110000111010011111010100000;
filter5[4][917] = 35'b00000001000101001000101001000100000;
filter5[4][918] = 35'b00000001101100010000110010000100000;
filter5[4][919] = 35'b11111110011111001110010101100100000;
filter5[4][920] = 35'b11111111101100100001110111110001100;
filter5[4][921] = 35'b00000000000001010010000100010010110;
filter5[4][922] = 35'b00000010101110011011011011000000000;
filter5[4][923] = 35'b00000000110110110111011010000110000;
filter5[4][924] = 35'b00000010001110100010111100011100000;
filter5[4][925] = 35'b00000000100000011100000101011011000;
filter5[4][926] = 35'b11111010110110101001000010010000000;
filter5[4][927] = 35'b11111100000101110100101001110000000;
filter5[4][928] = 35'b00000100111111101110011011101000000;
filter5[4][929] = 35'b11111111011000110001111111110000000;
filter5[4][930] = 35'b00000000111110110111110111010000000;
filter5[4][931] = 35'b11111111011101000001111011100010000;
filter5[4][932] = 35'b11111110000010011101011001111010000;
filter5[4][933] = 35'b00000000011111100100000011000101100;
filter5[4][934] = 35'b11111011110110001111000100110000000;
filter5[4][935] = 35'b11111000100110010001110001000000000;
filter5[4][936] = 35'b11111111100110011101101000011001100;
filter5[4][937] = 35'b00000011000101101010011101010100000;
filter5[4][938] = 35'b11111101101110111111101011001100000;
filter5[4][939] = 35'b00000011001110010010100110010100000;
filter5[4][940] = 35'b11111111011110110111101111000110000;
filter5[4][941] = 35'b11111101010111101011011011111100000;
filter5[4][942] = 35'b11111110010100000011001101011110000;
filter5[4][943] = 35'b11111001111101100001100110101000000;
filter5[4][944] = 35'b00000000100011001011101101101110000;
filter5[4][945] = 35'b00000001000011011000100010100100000;
filter5[4][946] = 35'b00000000000010110100011010110001101;
filter5[4][947] = 35'b00000000010011110010111010011000100;
filter5[4][948] = 35'b00000000100110101011001111010010000;
filter5[4][949] = 35'b11111100101110100101101111000000000;
filter5[4][950] = 35'b11111111101110110110111011111101100;
filter5[4][951] = 35'b11111111110011000000101101011000000;
filter5[4][952] = 35'b00000001000101011010110001101000000;
filter5[4][953] = 35'b00000111011000001110001001001000000;
filter5[4][954] = 35'b11111101100100111010000001111100000;
filter5[4][955] = 35'b11111111000001111100110001101100000;
filter5[4][956] = 35'b11111110110001001100101110011000000;
filter5[4][957] = 35'b00000001010010011100011011010110000;
filter5[4][958] = 35'b11111100000110000000100111101100000;
filter5[4][959] = 35'b11110100010110011111100101010000000;
filter5[4][960] = 35'b11111101010011010001110001011100000;
filter5[4][961] = 35'b00000001000011000011011111010110000;
filter5[4][962] = 35'b00001000010010100110001011000000000;
filter5[4][963] = 35'b00000110000010010001010100101000000;
filter5[4][964] = 35'b00000100010110001111101100000000000;
filter5[4][965] = 35'b11111100011100111111111000101100000;
filter5[4][966] = 35'b00000001010110110100100110111000000;
filter5[4][967] = 35'b11111011111011001000011001100000000;
filter5[4][968] = 35'b00000101110010110100011001101000000;
filter5[4][969] = 35'b00000011011101000100011111001000000;
filter5[4][970] = 35'b11111011100011101100000111100000000;
filter5[4][971] = 35'b11111100111111111011011100100100000;
filter5[4][972] = 35'b11111111001001110101001000111100000;
filter5[4][973] = 35'b00000011011010110000100000100100000;
filter5[4][974] = 35'b00000010100110001110010000001100000;
filter5[4][975] = 35'b11111110111000100111110000100000000;
filter5[4][976] = 35'b11111100100001011000001011011100000;
filter5[4][977] = 35'b11111110110010100000101011111110000;
filter5[4][978] = 35'b00000000111010110011011011011111000;
filter5[4][979] = 35'b11111111101110101011101010101001100;
filter5[4][980] = 35'b00000000001100111011000101001100100;
filter5[4][981] = 35'b11111110100010111110011111001110000;
filter5[4][982] = 35'b00000010111000011111011010110000000;
filter5[4][983] = 35'b11111100110101010111000101111000000;
filter5[4][984] = 35'b00000001011101110000010011011110000;
filter5[4][985] = 35'b11111110110110110001010011001110000;
filter5[4][986] = 35'b00000100000001001110010110100000000;
filter5[4][987] = 35'b11111110001011011001011011010100000;
filter5[4][988] = 35'b00000000100111100000101000000010000;
filter5[4][989] = 35'b00000010110111110000010000001100000;
filter5[4][990] = 35'b11111111110001010100000010100100000;
filter5[4][991] = 35'b00000000110110101110000101100101000;
filter5[4][992] = 35'b11111100111101011101111101110100000;
filter5[4][993] = 35'b11111111111110001011011010001111001;
filter5[4][994] = 35'b11111111000011110111100011010100000;
filter5[4][995] = 35'b00000011101100001100101111011100000;
filter5[4][996] = 35'b11111100101010101101110100110000000;
filter5[4][997] = 35'b11111000100010101111110110011000000;
filter5[4][998] = 35'b00000000010101101001000010011111100;
filter5[4][999] = 35'b11111101101100100010100011101100000;
filter5[4][1000] = 35'b11111110000010110010100000001000000;
filter5[4][1001] = 35'b00000100000000100000100011100000000;
filter5[4][1002] = 35'b00000001111101100001000000001010000;
filter5[4][1003] = 35'b11111111010000100101100111010100000;
filter5[4][1004] = 35'b00000010001111000110100110100000000;
filter5[4][1005] = 35'b11111011001111101000001111010000000;
filter5[4][1006] = 35'b11111011000000010000001000011000000;
filter5[4][1007] = 35'b11111011111111011010000110000000000;
filter5[4][1008] = 35'b11111100001011101011100010001000000;
filter5[4][1009] = 35'b00000101100000000001010010100000000;
filter5[4][1010] = 35'b00000011101001101011010001011100000;
filter5[4][1011] = 35'b11111111001100001110011110111000000;
filter5[4][1012] = 35'b00000010110110001110011100001000000;
filter5[4][1013] = 35'b11110111001110111000000000100000000;
filter5[4][1014] = 35'b11111110010100011111100010000010000;
filter5[4][1015] = 35'b11111010010000101110000000100000000;
filter5[4][1016] = 35'b11111010111110101111011101110000000;
filter5[4][1017] = 35'b00000001011110010101101001011110000;
filter5[4][1018] = 35'b00001000110010101101110000100000000;
filter5[4][1019] = 35'b11111011111010011001110010111000000;
filter5[4][1020] = 35'b00000001111011111011010101011100000;
filter5[4][1021] = 35'b11111111100001001101010010000000000;
filter5[4][1022] = 35'b11111001001101101110111001101000000;
filter5[4][1023] = 35'b11110101010100111001111000110000000;
filter5[5][0] = 35'b00000010010101111001111000101100000;
filter5[5][1] = 35'b00000001010101000100101101101110000;
filter5[5][2] = 35'b11111011100111000101010000101000000;
filter5[5][3] = 35'b11111010110101011110101110010000000;
filter5[5][4] = 35'b11111111111001011010100000001010010;
filter5[5][5] = 35'b00000010001101110000110111110000000;
filter5[5][6] = 35'b00000001111111000100110010101100000;
filter5[5][7] = 35'b00000110100100111010000000100000000;
filter5[5][8] = 35'b11111110011010111000000101000100000;
filter5[5][9] = 35'b00000001001010000010001011010000000;
filter5[5][10] = 35'b11111000010110001011100111110000000;
filter5[5][11] = 35'b11111111101011101000110111111110000;
filter5[5][12] = 35'b00000010111111100010100011000100000;
filter5[5][13] = 35'b00000110100000111010111010011000000;
filter5[5][14] = 35'b11111000000111110100001001100000000;
filter5[5][15] = 35'b00000110111110010000000111001000000;
filter5[5][16] = 35'b00000010001001101101100010010100000;
filter5[5][17] = 35'b00000000101010001100101100101010000;
filter5[5][18] = 35'b11111011100001110000001010110000000;
filter5[5][19] = 35'b11111110111100000111001010111000000;
filter5[5][20] = 35'b11111111010111101011000010101101000;
filter5[5][21] = 35'b00000010101110000100011010011000000;
filter5[5][22] = 35'b00000000011000100011011000001100100;
filter5[5][23] = 35'b11111110000101001010111110011110000;
filter5[5][24] = 35'b11111110010010100101011101010010000;
filter5[5][25] = 35'b11111110010010010111110001010110000;
filter5[5][26] = 35'b00000010011101010010111010111100000;
filter5[5][27] = 35'b00000001111111110100111111011100000;
filter5[5][28] = 35'b11111111100101100000000111100001000;
filter5[5][29] = 35'b11111111011011011001011111111110000;
filter5[5][30] = 35'b00000111111001101000110100000000000;
filter5[5][31] = 35'b00000101010111101010010000001000000;
filter5[5][32] = 35'b00000001010001110000110010111110000;
filter5[5][33] = 35'b11111110110000110000000110000110000;
filter5[5][34] = 35'b00000001001000011100000010001000000;
filter5[5][35] = 35'b11111111111011010100111011001000110;
filter5[5][36] = 35'b11111111100001101000000100011011100;
filter5[5][37] = 35'b11111101000111000000000101110100000;
filter5[5][38] = 35'b11111110000110110011011010101100000;
filter5[5][39] = 35'b00000010110010011001111100100100000;
filter5[5][40] = 35'b11111101111110011011011110010100000;
filter5[5][41] = 35'b11111110111010111111010110110100000;
filter5[5][42] = 35'b11111110100111100111100100001000000;
filter5[5][43] = 35'b11111111010011101101011101000111000;
filter5[5][44] = 35'b00000011011101101101010011101000000;
filter5[5][45] = 35'b11111111001111000010110100000001000;
filter5[5][46] = 35'b11111110001101010101101110101110000;
filter5[5][47] = 35'b00000100011011101100101000001000000;
filter5[5][48] = 35'b00000011000110010000001111000100000;
filter5[5][49] = 35'b00000010111000010101010110011000000;
filter5[5][50] = 35'b11111111110010110111100111111001000;
filter5[5][51] = 35'b11111111100101111010000011100111100;
filter5[5][52] = 35'b00000001000111010001111001100100000;
filter5[5][53] = 35'b11111000011011001010011001111000000;
filter5[5][54] = 35'b00000110001010100001100101101000000;
filter5[5][55] = 35'b00000011110001001110010111001000000;
filter5[5][56] = 35'b00000100010001001011111110011000000;
filter5[5][57] = 35'b00000001000001011101010111110000000;
filter5[5][58] = 35'b00000001010110101010010011111010000;
filter5[5][59] = 35'b11111100101100100100100011110100000;
filter5[5][60] = 35'b00000000001110100001100101101001010;
filter5[5][61] = 35'b00000111011110110011000000010000000;
filter5[5][62] = 35'b00000100111101000111110011011000000;
filter5[5][63] = 35'b00000110001100100001011111011000000;
filter5[5][64] = 35'b00000100100110111000111011000000000;
filter5[5][65] = 35'b00000000011110101001001001010110100;
filter5[5][66] = 35'b11111101100010100101010011010100000;
filter5[5][67] = 35'b11111101000110010101000001110000000;
filter5[5][68] = 35'b00000001000011001101011110011110000;
filter5[5][69] = 35'b00000001111011000110111011111000000;
filter5[5][70] = 35'b00000000010000011000011110011100100;
filter5[5][71] = 35'b00000101100111101011110010110000000;
filter5[5][72] = 35'b11111111011100011111011011001111000;
filter5[5][73] = 35'b11111100111011001010010001010100000;
filter5[5][74] = 35'b11111000011100011110010010100000000;
filter5[5][75] = 35'b11111110111001101011000000111110000;
filter5[5][76] = 35'b11111100100100101011100111100100000;
filter5[5][77] = 35'b00000010010010101111001000100100000;
filter5[5][78] = 35'b11111110111011101010100010001010000;
filter5[5][79] = 35'b00000011010000011010011111001000000;
filter5[5][80] = 35'b11111110011101111011011100111000000;
filter5[5][81] = 35'b11111111100100101010010011110010000;
filter5[5][82] = 35'b11111101100000011110110010010000000;
filter5[5][83] = 35'b11111111101010010101001100011100000;
filter5[5][84] = 35'b00000000011111100111111010001001000;
filter5[5][85] = 35'b00000001111000111010011001101110000;
filter5[5][86] = 35'b00000010000010101010001101110000000;
filter5[5][87] = 35'b11111100100000111001010011011100000;
filter5[5][88] = 35'b00000001000010001101101111100100000;
filter5[5][89] = 35'b11111011000001010011101101111000000;
filter5[5][90] = 35'b00000001100011101000100101101100000;
filter5[5][91] = 35'b11111111001101100111011111011101000;
filter5[5][92] = 35'b00000001010000101010110010111100000;
filter5[5][93] = 35'b00000011000011001010010001000000000;
filter5[5][94] = 35'b00000001110110000010010010101000000;
filter5[5][95] = 35'b11111111010110001011000011110001000;
filter5[5][96] = 35'b00000000010000001100101100110010000;
filter5[5][97] = 35'b11111101110001110010011010010000000;
filter5[5][98] = 35'b00000010111101100101001010100000000;
filter5[5][99] = 35'b11111110011000010001000111011100000;
filter5[5][100] = 35'b00000001001001000010101101100000000;
filter5[5][101] = 35'b11111110001110111011111110101110000;
filter5[5][102] = 35'b11111101111010111001001000110000000;
filter5[5][103] = 35'b11111100101011101101000110101000000;
filter5[5][104] = 35'b11111110011111000101110110010010000;
filter5[5][105] = 35'b11111101111110100011011000000000000;
filter5[5][106] = 35'b11111110010010011111001010011110000;
filter5[5][107] = 35'b11111101010011101111100000000000000;
filter5[5][108] = 35'b00000001100101110111110111010000000;
filter5[5][109] = 35'b11111111100111000101001010111100100;
filter5[5][110] = 35'b00000010110010001100110111111000000;
filter5[5][111] = 35'b00000011011110101010100110101000000;
filter5[5][112] = 35'b00000010000100101001010011100100000;
filter5[5][113] = 35'b11111110101100010100110011110110000;
filter5[5][114] = 35'b00000000001011000010010100011100100;
filter5[5][115] = 35'b11111101100010000001001110101000000;
filter5[5][116] = 35'b00000000110111010111001100001001000;
filter5[5][117] = 35'b00000000010010000011111111000101000;
filter5[5][118] = 35'b00000011101001011100110101000000000;
filter5[5][119] = 35'b00001000001101010111010111010000000;
filter5[5][120] = 35'b00000000110000010110110001111110000;
filter5[5][121] = 35'b11111111100110110100111111110000100;
filter5[5][122] = 35'b00000010110010010010010100000100000;
filter5[5][123] = 35'b11111011110000101000001101001000000;
filter5[5][124] = 35'b00000011000010111110110110011000000;
filter5[5][125] = 35'b11111101011100101000110011001100000;
filter5[5][126] = 35'b11111101100100000010101010011000000;
filter5[5][127] = 35'b00001000111100001101110001000000000;
filter5[5][128] = 35'b11111011101101000000111111001000000;
filter5[5][129] = 35'b11111110001101011101111000110010000;
filter5[5][130] = 35'b11110101111100001111011010110000000;
filter5[5][131] = 35'b11101011001100111100101111100000000;
filter5[5][132] = 35'b00000001011111001110110110100000000;
filter5[5][133] = 35'b00000011100111011000110001011000000;
filter5[5][134] = 35'b00000010111011000010011011001000000;
filter5[5][135] = 35'b00001001110100101110100110010000000;
filter5[5][136] = 35'b11111010011101011101010101011000000;
filter5[5][137] = 35'b11101001111110101000100111000000000;
filter5[5][138] = 35'b11101001111010101111011001100000000;
filter5[5][139] = 35'b11111110001011101111111111010100000;
filter5[5][140] = 35'b11111111011110101111010000101111000;
filter5[5][141] = 35'b00000011001100001011101110110000000;
filter5[5][142] = 35'b00000001111011100100111000110000000;
filter5[5][143] = 35'b11111100111000010000101100011100000;
filter5[5][144] = 35'b00000010100101100011100011000000000;
filter5[5][145] = 35'b11111100100001110010101100010000000;
filter5[5][146] = 35'b11111011000101000101110001110000000;
filter5[5][147] = 35'b00000010110101101100001010110100000;
filter5[5][148] = 35'b00000000100010110010111010010101000;
filter5[5][149] = 35'b00000011110011000000001110000000000;
filter5[5][150] = 35'b11111110010011110100011010000100000;
filter5[5][151] = 35'b00000000000110110001100001110010001;
filter5[5][152] = 35'b11111100011000111010011100110100000;
filter5[5][153] = 35'b11110111110001101010111001000000000;
filter5[5][154] = 35'b00000000110100100111110110011111000;
filter5[5][155] = 35'b00000100000011011101000100000000000;
filter5[5][156] = 35'b00000000010101100001011011011010000;
filter5[5][157] = 35'b00000000001111000111001110010010000;
filter5[5][158] = 35'b11111111000011000100000110000111000;
filter5[5][159] = 35'b00000001010000101010101011001000000;
filter5[5][160] = 35'b00000001010001110000010010000010000;
filter5[5][161] = 35'b11111100001110010000100001111100000;
filter5[5][162] = 35'b00000001001001000111010111010010000;
filter5[5][163] = 35'b11110110110101011111110011110000000;
filter5[5][164] = 35'b00000001001010010110101111111110000;
filter5[5][165] = 35'b11111011101101111000000011001000000;
filter5[5][166] = 35'b11111110011011111100111010101110000;
filter5[5][167] = 35'b11110110001000011110000111000000000;
filter5[5][168] = 35'b11111010101100100101100110110000000;
filter5[5][169] = 35'b00000110110001111011101101011000000;
filter5[5][170] = 35'b11111101100010111111110001010000000;
filter5[5][171] = 35'b11111000001111010001011011100000000;
filter5[5][172] = 35'b11111001111101000011000101101000000;
filter5[5][173] = 35'b00000110011100101000100111000000000;
filter5[5][174] = 35'b00000110000100001011011010110000000;
filter5[5][175] = 35'b00000110001110011001111000111000000;
filter5[5][176] = 35'b11111100101001010110000100100100000;
filter5[5][177] = 35'b11111111101110011001100010100111100;
filter5[5][178] = 35'b11111011100100000100010011010000000;
filter5[5][179] = 35'b11110100100111101110111000110000000;
filter5[5][180] = 35'b11010111000101100001001100000000000;
filter5[5][181] = 35'b00000010100011010110001001101100000;
filter5[5][182] = 35'b00001000001101111110001000100000000;
filter5[5][183] = 35'b11111101101100010001100001010100000;
filter5[5][184] = 35'b11111001101000110110100111101000000;
filter5[5][185] = 35'b11111111100101111111101011111111000;
filter5[5][186] = 35'b11111111001000001100100000011101000;
filter5[5][187] = 35'b11111100010100100111001100001100000;
filter5[5][188] = 35'b00000100101101011000001001000000000;
filter5[5][189] = 35'b11110100101111101010001111100000000;
filter5[5][190] = 35'b00010001000011100101010011000000000;
filter5[5][191] = 35'b00001110010100000100000011010000000;
filter5[5][192] = 35'b11111111001011000000001000110101000;
filter5[5][193] = 35'b00000001110000111111010100001000000;
filter5[5][194] = 35'b11110010100010100010111000010000000;
filter5[5][195] = 35'b11111000001011101000000000100000000;
filter5[5][196] = 35'b11110100111100101100010011010000000;
filter5[5][197] = 35'b00000010000100110001011011000000000;
filter5[5][198] = 35'b00000110111000001110110001001000000;
filter5[5][199] = 35'b00000100100110111110101100110000000;
filter5[5][200] = 35'b00000000001000110000101011101110100;
filter5[5][201] = 35'b00000011111111110110101010110100000;
filter5[5][202] = 35'b11110001100011011111111001000000000;
filter5[5][203] = 35'b11111000100110110001100100000000000;
filter5[5][204] = 35'b00000000110101001001010101010111000;
filter5[5][205] = 35'b00000100001101011001100100011000000;
filter5[5][206] = 35'b00000001010001110110011111001000000;
filter5[5][207] = 35'b11111001000001100010000010101000000;
filter5[5][208] = 35'b11111001010001001010001001110000000;
filter5[5][209] = 35'b11111001000110011010110101101000000;
filter5[5][210] = 35'b11111101000101000110111011001100000;
filter5[5][211] = 35'b11111110101011101100110100000010000;
filter5[5][212] = 35'b11111011011111010001111101011000000;
filter5[5][213] = 35'b00001001010111000111000011100000000;
filter5[5][214] = 35'b00000011010100011001101110110000000;
filter5[5][215] = 35'b11111110011101011000010100010010000;
filter5[5][216] = 35'b11111010100001001010001110110000000;
filter5[5][217] = 35'b11111101001101000000111110011100000;
filter5[5][218] = 35'b11111100011111011101000001110000000;
filter5[5][219] = 35'b00000001000000000001110000100110000;
filter5[5][220] = 35'b11111111001011011101111101100000000;
filter5[5][221] = 35'b11111101100000110011110110100100000;
filter5[5][222] = 35'b00000000011011110110101010011100100;
filter5[5][223] = 35'b11111110111110101100011001100100000;
filter5[5][224] = 35'b11110111110100011011100101100000000;
filter5[5][225] = 35'b11111111110101100000010100010000110;
filter5[5][226] = 35'b11111100111010001110110001111100000;
filter5[5][227] = 35'b00000001101101011011100010100010000;
filter5[5][228] = 35'b11111110110100001100111000111010000;
filter5[5][229] = 35'b00000000111011101010000011000111000;
filter5[5][230] = 35'b00000000110100101001011100101000000;
filter5[5][231] = 35'b00000011100010100000101010000000000;
filter5[5][232] = 35'b11101110111000011100111111100000000;
filter5[5][233] = 35'b11111110011100111000100111111100000;
filter5[5][234] = 35'b11111101110000011000001101111100000;
filter5[5][235] = 35'b11111111110111100010101100101100010;
filter5[5][236] = 35'b00000001010110100000010100110010000;
filter5[5][237] = 35'b00000011000100101111000110100000000;
filter5[5][238] = 35'b11111011010101001110010111000000000;
filter5[5][239] = 35'b00000000110110101101100100101011000;
filter5[5][240] = 35'b11111001111010110111110110101000000;
filter5[5][241] = 35'b00000001011101100111010110000010000;
filter5[5][242] = 35'b11111100011010001001010101100000000;
filter5[5][243] = 35'b11111101111000100010000101100000000;
filter5[5][244] = 35'b11111111010101011111100001101101000;
filter5[5][245] = 35'b00000001011110100111111001110010000;
filter5[5][246] = 35'b00000010110111111110010000100100000;
filter5[5][247] = 35'b00000001101111101111101011000110000;
filter5[5][248] = 35'b11111010110001001111101101010000000;
filter5[5][249] = 35'b11111010001101001011000101100000000;
filter5[5][250] = 35'b00000010011111111000001000110100000;
filter5[5][251] = 35'b00000011000100100110010011000100000;
filter5[5][252] = 35'b11111100010100100101010000101000000;
filter5[5][253] = 35'b00000010001110010001111110001000000;
filter5[5][254] = 35'b11111111001010010011001101000001000;
filter5[5][255] = 35'b00000011101010011001101110000100000;
filter5[5][256] = 35'b00000001100011100010010100010100000;
filter5[5][257] = 35'b11111111001010000010000010001001000;
filter5[5][258] = 35'b11111110000111100010111011000110000;
filter5[5][259] = 35'b11110101111110001101110001010000000;
filter5[5][260] = 35'b11110110010111011001111010110000000;
filter5[5][261] = 35'b00001000100111101000010110100000000;
filter5[5][262] = 35'b00000111110001001100110010010000000;
filter5[5][263] = 35'b00000001001000111110011000110100000;
filter5[5][264] = 35'b11111110110100101000001010001110000;
filter5[5][265] = 35'b11111100000110000100010011011000000;
filter5[5][266] = 35'b11110110100001111110111111110000000;
filter5[5][267] = 35'b00000001000001101010100001000010000;
filter5[5][268] = 35'b00000110101100000001101111000000000;
filter5[5][269] = 35'b00000010010011100010000011101100000;
filter5[5][270] = 35'b11111010111010110101000010011000000;
filter5[5][271] = 35'b11111100101010100100001100011000000;
filter5[5][272] = 35'b11111000111010100100010110100000000;
filter5[5][273] = 35'b11111001111011110101100000001000000;
filter5[5][274] = 35'b11111110000100111110111001011000000;
filter5[5][275] = 35'b11111101011111101110001011010100000;
filter5[5][276] = 35'b00000001100011010110000110101010000;
filter5[5][277] = 35'b00000010011111000010000111111100000;
filter5[5][278] = 35'b11111110001110100010110111111110000;
filter5[5][279] = 35'b11110010100110000010010110100000000;
filter5[5][280] = 35'b11110111001000100001101001000000000;
filter5[5][281] = 35'b11111010100011100100011001001000000;
filter5[5][282] = 35'b00000100010011011101001001110000000;
filter5[5][283] = 35'b00000010010101111011010110110000000;
filter5[5][284] = 35'b11111111000100000111010110110001000;
filter5[5][285] = 35'b11111110100000011100000010101100000;
filter5[5][286] = 35'b11111011010010110111011011101000000;
filter5[5][287] = 35'b00000000101001111100001011111010000;
filter5[5][288] = 35'b11110011111110011000011001010000000;
filter5[5][289] = 35'b00000000000110111110010111100111000;
filter5[5][290] = 35'b00000000011001001111101101011101100;
filter5[5][291] = 35'b00000011000011010001101001100000000;
filter5[5][292] = 35'b11111111010011110101100110111000000;
filter5[5][293] = 35'b00000001000111011000000101111100000;
filter5[5][294] = 35'b11111111100010101000110010101111000;
filter5[5][295] = 35'b00000100001001111010100110011000000;
filter5[5][296] = 35'b11101111010011100001111101000000000;
filter5[5][297] = 35'b11110111110111110001000011000000000;
filter5[5][298] = 35'b11111011010001100000100001001000000;
filter5[5][299] = 35'b11111111000110000001111000110011000;
filter5[5][300] = 35'b00000001110111100001011011111110000;
filter5[5][301] = 35'b00000011001011001000111111011100000;
filter5[5][302] = 35'b00000001000000011111101101101100000;
filter5[5][303] = 35'b00000011011110101110011100100000000;
filter5[5][304] = 35'b11111101001100010001110110011100000;
filter5[5][305] = 35'b11111110001100001100101111001110000;
filter5[5][306] = 35'b11111110110011110111001110100100000;
filter5[5][307] = 35'b11111100101010110100111100011000000;
filter5[5][308] = 35'b00000001011000101110111110000010000;
filter5[5][309] = 35'b00000010111010111011011000111000000;
filter5[5][310] = 35'b00000000000011000111100011000100100;
filter5[5][311] = 35'b00000101000011001000101101000000000;
filter5[5][312] = 35'b11110110001000010100101100110000000;
filter5[5][313] = 35'b11111000000100011001011000011000000;
filter5[5][314] = 35'b00000101011101011101110010101000000;
filter5[5][315] = 35'b11111100101001111100000100010100000;
filter5[5][316] = 35'b11111100101100111101000010110000000;
filter5[5][317] = 35'b11111010110111110111001111101000000;
filter5[5][318] = 35'b11111110000000010011000111101100000;
filter5[5][319] = 35'b00000100011001010001101100100000000;
filter5[5][320] = 35'b00000100011001001100000110100000000;
filter5[5][321] = 35'b00000001101011110110110101100110000;
filter5[5][322] = 35'b11111010100010011011101011110000000;
filter5[5][323] = 35'b00000000010001110010010101110001000;
filter5[5][324] = 35'b00000001100100111101101100100000000;
filter5[5][325] = 35'b00000010110000111111101010000100000;
filter5[5][326] = 35'b00000000000111010111000000100001000;
filter5[5][327] = 35'b00000111100000100111111100110000000;
filter5[5][328] = 35'b11111111100110001111000101001111000;
filter5[5][329] = 35'b11111110010010000101101111101100000;
filter5[5][330] = 35'b11110111101110011101111101110000000;
filter5[5][331] = 35'b11111001100101001001100001110000000;
filter5[5][332] = 35'b11111110011000011000111110110100000;
filter5[5][333] = 35'b00000010011001001110110111011000000;
filter5[5][334] = 35'b00000000011010010111111100100100000;
filter5[5][335] = 35'b11111110100101111100010011110010000;
filter5[5][336] = 35'b00000010001011000000000011011000000;
filter5[5][337] = 35'b00000001010001101010111101101000000;
filter5[5][338] = 35'b11111110111001111111001000001100000;
filter5[5][339] = 35'b11111111010101100101100111111001000;
filter5[5][340] = 35'b11111111101101011110100010011011000;
filter5[5][341] = 35'b00000101011011111011110100001000000;
filter5[5][342] = 35'b11111111101111010001000100111111000;
filter5[5][343] = 35'b11111101000101000101001000101100000;
filter5[5][344] = 35'b00000001110110010011001101001110000;
filter5[5][345] = 35'b11111111100101100011111101111001000;
filter5[5][346] = 35'b11111101100101010011000101111000000;
filter5[5][347] = 35'b00000100011110000111101110000000000;
filter5[5][348] = 35'b11111110100000101100000100110010000;
filter5[5][349] = 35'b00000010001101111010111011001100000;
filter5[5][350] = 35'b00000010001111111000010111000100000;
filter5[5][351] = 35'b11111110001110001000110000101110000;
filter5[5][352] = 35'b00000001110100101010111010011000000;
filter5[5][353] = 35'b11111111011000000001110011111101000;
filter5[5][354] = 35'b11111101000100111110100100101100000;
filter5[5][355] = 35'b11111111000101011000110100110110000;
filter5[5][356] = 35'b11111110110000011000000110011100000;
filter5[5][357] = 35'b00000000111000001100000100100011000;
filter5[5][358] = 35'b11111101110111100001101000010000000;
filter5[5][359] = 35'b00000000101110000010101000010001000;
filter5[5][360] = 35'b00000011011100010101001010100100000;
filter5[5][361] = 35'b11111111101001011001001101001011100;
filter5[5][362] = 35'b11111100001111001110001101101100000;
filter5[5][363] = 35'b11111111110100011100010111100001100;
filter5[5][364] = 35'b00000001000001111010101101100000000;
filter5[5][365] = 35'b00000001001100000101101110100010000;
filter5[5][366] = 35'b11111110100000101101111101010110000;
filter5[5][367] = 35'b00000010101111010000010111010100000;
filter5[5][368] = 35'b00000000010101101111000101010101100;
filter5[5][369] = 35'b00000000001101101110100111011011100;
filter5[5][370] = 35'b00000000011100001011011111110011000;
filter5[5][371] = 35'b11111110011101110100000001100000000;
filter5[5][372] = 35'b00000000010100001000011111010011100;
filter5[5][373] = 35'b11111100111100000100110011101100000;
filter5[5][374] = 35'b00000100001000011110001111001000000;
filter5[5][375] = 35'b00000011100010100110111010001000000;
filter5[5][376] = 35'b11111110111010101100011010010110000;
filter5[5][377] = 35'b11111101101011100000111000100000000;
filter5[5][378] = 35'b00000011010100110010101011100100000;
filter5[5][379] = 35'b00000000010111101111011010010100100;
filter5[5][380] = 35'b11111111000011111011100011001001000;
filter5[5][381] = 35'b00000100111101110100001111000000000;
filter5[5][382] = 35'b11111111101010011001000001000010000;
filter5[5][383] = 35'b00000101000010011110101100111000000;
filter5[5][384] = 35'b00000000100100001101111110000001000;
filter5[5][385] = 35'b00000010000101101001010111000100000;
filter5[5][386] = 35'b00000000001111000011110101011110100;
filter5[5][387] = 35'b00000011010110101111111101110100000;
filter5[5][388] = 35'b00000011101000000110100111011100000;
filter5[5][389] = 35'b00000001010001101110101010000010000;
filter5[5][390] = 35'b00000000100110101101011000110010000;
filter5[5][391] = 35'b00000000011101110111011000011100100;
filter5[5][392] = 35'b00000000101111111000000000111110000;
filter5[5][393] = 35'b00000010010000111011010001010000000;
filter5[5][394] = 35'b00000000001000000111101000111110010;
filter5[5][395] = 35'b00000010110011011010110010001100000;
filter5[5][396] = 35'b00000001000010001111111010110100000;
filter5[5][397] = 35'b11111110000111111010001110110010000;
filter5[5][398] = 35'b00000000111110111111111000010111000;
filter5[5][399] = 35'b11111111000001011000010111101100000;
filter5[5][400] = 35'b11111110001001011111100111101110000;
filter5[5][401] = 35'b11111111001101101111110111011111000;
filter5[5][402] = 35'b00000001001000110010111111100000000;
filter5[5][403] = 35'b00000001001010010110001110101000000;
filter5[5][404] = 35'b11111110010110110011100111010010000;
filter5[5][405] = 35'b11111100000110000100000010111000000;
filter5[5][406] = 35'b11111111110000000100011111001001010;
filter5[5][407] = 35'b11111100101010011111111111101100000;
filter5[5][408] = 35'b11111111100110001111110101110011000;
filter5[5][409] = 35'b11111111000001001111001110010110000;
filter5[5][410] = 35'b11111011111111010011011101011000000;
filter5[5][411] = 35'b11111101110100000110100011011000000;
filter5[5][412] = 35'b00000010000100101110110010111100000;
filter5[5][413] = 35'b11111111111000111010001000110000011;
filter5[5][414] = 35'b11111111101110101011101011001010000;
filter5[5][415] = 35'b11111101110001111101011101101000000;
filter5[5][416] = 35'b11111101100110011101101100100100000;
filter5[5][417] = 35'b00000010001010111000111100010100000;
filter5[5][418] = 35'b00000000101111011101001001101010000;
filter5[5][419] = 35'b11111111101011010011011100010011100;
filter5[5][420] = 35'b00000000000100001010010111101101111;
filter5[5][421] = 35'b11111100000100110101001101110000000;
filter5[5][422] = 35'b11110110010110000011010000010000000;
filter5[5][423] = 35'b11111011101000101001100101111000000;
filter5[5][424] = 35'b00000001110011000101101111000000000;
filter5[5][425] = 35'b00000010000111111001011010000100000;
filter5[5][426] = 35'b11111111010111110100101111010000000;
filter5[5][427] = 35'b00000000000100111111011101011100100;
filter5[5][428] = 35'b11111010101000111001010100101000000;
filter5[5][429] = 35'b11111000111100000110001101100000000;
filter5[5][430] = 35'b11111100100100101111000111011100000;
filter5[5][431] = 35'b00000011001110010100000100011000000;
filter5[5][432] = 35'b00000001010000010001100101000010000;
filter5[5][433] = 35'b00000000011010100011001100110101000;
filter5[5][434] = 35'b00000010101111100101000101010100000;
filter5[5][435] = 35'b00000010001011001110101011011100000;
filter5[5][436] = 35'b11111110011101111101011110110100000;
filter5[5][437] = 35'b11111100110100111011100110011000000;
filter5[5][438] = 35'b11111101111010111111010001100100000;
filter5[5][439] = 35'b00000100000110100000100111111000000;
filter5[5][440] = 35'b00000010100000111001101011010000000;
filter5[5][441] = 35'b00000001001100001100110000110000000;
filter5[5][442] = 35'b11111101111100010011101111001000000;
filter5[5][443] = 35'b00000110011110111000011001000000000;
filter5[5][444] = 35'b00000000100111101101110011011101000;
filter5[5][445] = 35'b00000100111101111111100110001000000;
filter5[5][446] = 35'b00000010100001111000111000100100000;
filter5[5][447] = 35'b00000111011001000010101100100000000;
filter5[5][448] = 35'b11111110110011001000010001010100000;
filter5[5][449] = 35'b00000101000101010001110101001000000;
filter5[5][450] = 35'b11111010010101011101001000101000000;
filter5[5][451] = 35'b11111101101101001000001011011000000;
filter5[5][452] = 35'b11111100010001001011110110101100000;
filter5[5][453] = 35'b11111100001001101011001001000100000;
filter5[5][454] = 35'b11111111111110111010000110111111010;
filter5[5][455] = 35'b11111101101100110001011010011100000;
filter5[5][456] = 35'b00000101100100000101101010010000000;
filter5[5][457] = 35'b00000000110001000110000100110011000;
filter5[5][458] = 35'b00000101110010110101101001010000000;
filter5[5][459] = 35'b00000110110100000000110111000000000;
filter5[5][460] = 35'b11111111011011010110000101001110000;
filter5[5][461] = 35'b00000101001110000110100000101000000;
filter5[5][462] = 35'b00000100011011001001000000110000000;
filter5[5][463] = 35'b11111110100100110010011101010110000;
filter5[5][464] = 35'b11111101010111100001101010100000000;
filter5[5][465] = 35'b11111101001010101011100000111100000;
filter5[5][466] = 35'b00000001100100110100010100011000000;
filter5[5][467] = 35'b00000111000100111011000100110000000;
filter5[5][468] = 35'b11111010001100111010000001001000000;
filter5[5][469] = 35'b00001001101011001001111111100000000;
filter5[5][470] = 35'b11110100010000001110111011010000000;
filter5[5][471] = 35'b00000100101000101110000111100000000;
filter5[5][472] = 35'b11111101000010000001011100011000000;
filter5[5][473] = 35'b00000101110110010010100011110000000;
filter5[5][474] = 35'b11111100110101000001010001111100000;
filter5[5][475] = 35'b11110110111111001101011011100000000;
filter5[5][476] = 35'b11110100111110010100101010100000000;
filter5[5][477] = 35'b11111111001101000101101110111001000;
filter5[5][478] = 35'b11110111100011011100010010000000000;
filter5[5][479] = 35'b11111010010010101000000010101000000;
filter5[5][480] = 35'b00000000011000010110001100101011100;
filter5[5][481] = 35'b11111111000011100110110110111000000;
filter5[5][482] = 35'b00000001111011011000111111010000000;
filter5[5][483] = 35'b11111100110111010101100000100100000;
filter5[5][484] = 35'b11110011111000001101110000010000000;
filter5[5][485] = 35'b11110101111101110100011101100000000;
filter5[5][486] = 35'b11111011010101101111101000100000000;
filter5[5][487] = 35'b00000001000000100111101000001100000;
filter5[5][488] = 35'b00000110100111000110000111100000000;
filter5[5][489] = 35'b11111101101101100101111001000000000;
filter5[5][490] = 35'b00000011011000000101101100100000000;
filter5[5][491] = 35'b00000110000011000100110001001000000;
filter5[5][492] = 35'b11111011011010110110111010010000000;
filter5[5][493] = 35'b11111111110110111101111100100001110;
filter5[5][494] = 35'b11111110111011110010000011001110000;
filter5[5][495] = 35'b00000100100000111111101111010000000;
filter5[5][496] = 35'b11111111100000001010110111011110000;
filter5[5][497] = 35'b11111101011001111111010110010100000;
filter5[5][498] = 35'b11111100001110100111110111100100000;
filter5[5][499] = 35'b11111101101000011011100011001000000;
filter5[5][500] = 35'b00000000101010111101101100010001000;
filter5[5][501] = 35'b00000010010000101100011101011000000;
filter5[5][502] = 35'b00000001000000110001010001000100000;
filter5[5][503] = 35'b00000010101110101100000000011000000;
filter5[5][504] = 35'b11111101001001001101001001101000000;
filter5[5][505] = 35'b00000000110010001010011001001001000;
filter5[5][506] = 35'b11111001010111110101111110100000000;
filter5[5][507] = 35'b00000001001100011101110110111010000;
filter5[5][508] = 35'b00000001100110000001011001100010000;
filter5[5][509] = 35'b00000011100011100001001000011100000;
filter5[5][510] = 35'b11111011011100101111111111001000000;
filter5[5][511] = 35'b00000010101110011101010100101000000;
filter5[5][512] = 35'b11111100011110101010000111100000000;
filter5[5][513] = 35'b00000100001110110101100101001000000;
filter5[5][514] = 35'b11111110101110000111000000101100000;
filter5[5][515] = 35'b11111110100010100000011010100110000;
filter5[5][516] = 35'b00000011110100101011001011010100000;
filter5[5][517] = 35'b00000100101010001010011101011000000;
filter5[5][518] = 35'b11111100110110000111101011110000000;
filter5[5][519] = 35'b11111110110101001110111100100110000;
filter5[5][520] = 35'b00000000100010100100100000000001000;
filter5[5][521] = 35'b00000001101100100001101101011100000;
filter5[5][522] = 35'b11111100001000100100010011010000000;
filter5[5][523] = 35'b11111100001101110111101111010000000;
filter5[5][524] = 35'b11111101001111010011100100101100000;
filter5[5][525] = 35'b00000000001001111101111101001001000;
filter5[5][526] = 35'b00000101100100100101110101100000000;
filter5[5][527] = 35'b11111110110110111110000011111000000;
filter5[5][528] = 35'b11111110101000000011010111100100000;
filter5[5][529] = 35'b00000001011100011110100010001000000;
filter5[5][530] = 35'b00000000010000110111110000011001000;
filter5[5][531] = 35'b11111110010110100010100111100110000;
filter5[5][532] = 35'b11111100111101011110111100110000000;
filter5[5][533] = 35'b11111100110110111011101010110100000;
filter5[5][534] = 35'b00000001111101100111000101001110000;
filter5[5][535] = 35'b00000010101001111110101101101100000;
filter5[5][536] = 35'b00000001110011110100010010101000000;
filter5[5][537] = 35'b11111011111110000111101111110000000;
filter5[5][538] = 35'b11111100010101000001111100101100000;
filter5[5][539] = 35'b11111100111011111010010101100100000;
filter5[5][540] = 35'b11111110000100000111101111101000000;
filter5[5][541] = 35'b00000010111110010110001111001100000;
filter5[5][542] = 35'b11111111000110100001011010110000000;
filter5[5][543] = 35'b00000011011100000111101010001000000;
filter5[5][544] = 35'b00000010100100011101000001011100000;
filter5[5][545] = 35'b00000001110101000000101100010010000;
filter5[5][546] = 35'b11111100011000101111101101000000000;
filter5[5][547] = 35'b11111111011100101000001000110100000;
filter5[5][548] = 35'b11111110001011001001000111111000000;
filter5[5][549] = 35'b11111111101101100011011010000111000;
filter5[5][550] = 35'b11111101000101111011100010111100000;
filter5[5][551] = 35'b11111111111101111110100000110010110;
filter5[5][552] = 35'b00000011110010010100011001000000000;
filter5[5][553] = 35'b00000000110010000110110110000011000;
filter5[5][554] = 35'b11111110100010111000101000101000000;
filter5[5][555] = 35'b11111011101010100001011011010000000;
filter5[5][556] = 35'b11111100000111000111100100000100000;
filter5[5][557] = 35'b11111111100110011010111010110010100;
filter5[5][558] = 35'b00000010010000100000010000100100000;
filter5[5][559] = 35'b00000100100111111001110000100000000;
filter5[5][560] = 35'b11111111001000100010011010011000000;
filter5[5][561] = 35'b00000010101011010001001011110100000;
filter5[5][562] = 35'b11111101011110001101001101010100000;
filter5[5][563] = 35'b11111111010011100001110100011000000;
filter5[5][564] = 35'b11111110110001001111111011000110000;
filter5[5][565] = 35'b00000010011110010011010110110000000;
filter5[5][566] = 35'b00000010011111111111011000010100000;
filter5[5][567] = 35'b00000010101011101010100000010100000;
filter5[5][568] = 35'b11111111001101010100110110000000000;
filter5[5][569] = 35'b00000010000100001010110010000000000;
filter5[5][570] = 35'b00000101111100010100001111010000000;
filter5[5][571] = 35'b11111101111101001011111101100100000;
filter5[5][572] = 35'b00000100111101010110010000101000000;
filter5[5][573] = 35'b00000001100101111011010001110100000;
filter5[5][574] = 35'b00000000110011110001110111101011000;
filter5[5][575] = 35'b00001010110101101011101011100000000;
filter5[5][576] = 35'b11111100011001110111110111011100000;
filter5[5][577] = 35'b00000001101010011000100100010000000;
filter5[5][578] = 35'b11111110011101111101000000101010000;
filter5[5][579] = 35'b11111111001110101101100110011111000;
filter5[5][580] = 35'b00000101000100100101001110110000000;
filter5[5][581] = 35'b00000011110011110111111110100100000;
filter5[5][582] = 35'b11111010010000110100011001000000000;
filter5[5][583] = 35'b11111011001100100001110010000000000;
filter5[5][584] = 35'b11111111111111001111100110011010111;
filter5[5][585] = 35'b00000000111111010000000000111001000;
filter5[5][586] = 35'b11111001010100100000111010000000000;
filter5[5][587] = 35'b11111011010011110110010110000000000;
filter5[5][588] = 35'b11111100110001001000100111101100000;
filter5[5][589] = 35'b00000000100100111011010111000111000;
filter5[5][590] = 35'b11111111101100001010101001001010100;
filter5[5][591] = 35'b00000000001110011010110011111100010;
filter5[5][592] = 35'b11111011000110101110011001011000000;
filter5[5][593] = 35'b11111101011111000001000111011000000;
filter5[5][594] = 35'b11111110101001101100111010010110000;
filter5[5][595] = 35'b11111100000000100100100110011000000;
filter5[5][596] = 35'b11111100100011000001000101001000000;
filter5[5][597] = 35'b11111111101011100110000101010011100;
filter5[5][598] = 35'b00000001000000001001001000111010000;
filter5[5][599] = 35'b00000001100000101001110111001110000;
filter5[5][600] = 35'b00000000011100111001111101000100000;
filter5[5][601] = 35'b11111111111011011110110100100001100;
filter5[5][602] = 35'b11111101010110100101111110010000000;
filter5[5][603] = 35'b00000001000001011100010001111000000;
filter5[5][604] = 35'b11111010111010001110010100000000000;
filter5[5][605] = 35'b00000000010010111101101011010001100;
filter5[5][606] = 35'b00000000111111010011101000111100000;
filter5[5][607] = 35'b11111111101111100111000010011111000;
filter5[5][608] = 35'b11111010111111001011011101111000000;
filter5[5][609] = 35'b11111100111000001100100101110000000;
filter5[5][610] = 35'b11111000011100000000101111010000000;
filter5[5][611] = 35'b00000000101101010011101101011111000;
filter5[5][612] = 35'b11111110111011001100000110001100000;
filter5[5][613] = 35'b00000010011001010100110110010000000;
filter5[5][614] = 35'b11111111010101100100001101101111000;
filter5[5][615] = 35'b00000011001011100010000111011100000;
filter5[5][616] = 35'b00000110100011001110100011111000000;
filter5[5][617] = 35'b11111101001011011001111001100100000;
filter5[5][618] = 35'b11111100111100000001110100001000000;
filter5[5][619] = 35'b00000001000110000001101110001100000;
filter5[5][620] = 35'b00000011000001111101011001110100000;
filter5[5][621] = 35'b11111111111010111011001000010010110;
filter5[5][622] = 35'b11111110111110001011011001001110000;
filter5[5][623] = 35'b00000010010011111000001100111100000;
filter5[5][624] = 35'b11111100010101101111110110101100000;
filter5[5][625] = 35'b11111010010110001101110000100000000;
filter5[5][626] = 35'b11111000111111011100110000101000000;
filter5[5][627] = 35'b11111110010100000010101110011010000;
filter5[5][628] = 35'b11111110100000101100011111101100000;
filter5[5][629] = 35'b00000011010011011000010001001000000;
filter5[5][630] = 35'b00000100010001010100111000001000000;
filter5[5][631] = 35'b00000001011010111101101110111100000;
filter5[5][632] = 35'b11111111101011111111001000100001100;
filter5[5][633] = 35'b11110111011010011101010101010000000;
filter5[5][634] = 35'b11111000100110101011010000001000000;
filter5[5][635] = 35'b00000101101010001101110010100000000;
filter5[5][636] = 35'b11111101101001100100111010011000000;
filter5[5][637] = 35'b00000001110001000000000001100100000;
filter5[5][638] = 35'b11111101000000010001101100011000000;
filter5[5][639] = 35'b00000100010101111110100100101000000;
filter5[5][640] = 35'b00000001111100100101111110101110000;
filter5[5][641] = 35'b00000011100101110110001110110100000;
filter5[5][642] = 35'b11111011001111001101011010001000000;
filter5[5][643] = 35'b00000101010011010010010110111000000;
filter5[5][644] = 35'b11111111001010100011001100001001000;
filter5[5][645] = 35'b11111011110000101000011000101000000;
filter5[5][646] = 35'b11111111111000100010110011001100010;
filter5[5][647] = 35'b00000100100001001011011111001000000;
filter5[5][648] = 35'b00000011010010011110110111011000000;
filter5[5][649] = 35'b00000010111010001010011100101000000;
filter5[5][650] = 35'b11111011011100001011100011110000000;
filter5[5][651] = 35'b00000100110001010101010101101000000;
filter5[5][652] = 35'b11111001100010111000011111101000000;
filter5[5][653] = 35'b11111100010011001010110010001000000;
filter5[5][654] = 35'b00000010111001100111101110110100000;
filter5[5][655] = 35'b11111000101110001111010011101000000;
filter5[5][656] = 35'b00000000111011001000100110100110000;
filter5[5][657] = 35'b00000010001110011101001110100000000;
filter5[5][658] = 35'b11111110101101011000010110001100000;
filter5[5][659] = 35'b11111111111010110110011000001010110;
filter5[5][660] = 35'b11111110100001101011011110100000000;
filter5[5][661] = 35'b11111110010010000100001101010110000;
filter5[5][662] = 35'b11111110000101101000000110000100000;
filter5[5][663] = 35'b00000100101011001110100001110000000;
filter5[5][664] = 35'b11111111010011100100110101001000000;
filter5[5][665] = 35'b00000000011000010111000011110000100;
filter5[5][666] = 35'b00000001001001010100011110111010000;
filter5[5][667] = 35'b11111111100001000010101111101000000;
filter5[5][668] = 35'b00000000010000001101011111111001100;
filter5[5][669] = 35'b11111111101100110111011000100011000;
filter5[5][670] = 35'b11111111001111110011000101100110000;
filter5[5][671] = 35'b11111110000010010010011010110110000;
filter5[5][672] = 35'b00000010011101010101101001001000000;
filter5[5][673] = 35'b00000011110001000111110000000000000;
filter5[5][674] = 35'b00000100110111101100001001110000000;
filter5[5][675] = 35'b11111101101000000000000010011100000;
filter5[5][676] = 35'b11111001010011000011001011010000000;
filter5[5][677] = 35'b00000000001111011101100010001101110;
filter5[5][678] = 35'b11111001100110110111111001010000000;
filter5[5][679] = 35'b00000000101010100011001010100111000;
filter5[5][680] = 35'b00000010010010001101100011111100000;
filter5[5][681] = 35'b00000001110001111001100000000010000;
filter5[5][682] = 35'b00000001011000001110011000010110000;
filter5[5][683] = 35'b00000000100010111110000010011111000;
filter5[5][684] = 35'b11111010100001000001111101110000000;
filter5[5][685] = 35'b11111100101001011001011110001100000;
filter5[5][686] = 35'b11111100000100111100110010100100000;
filter5[5][687] = 35'b00000010111011001110011111010100000;
filter5[5][688] = 35'b00000001110110011011000010111100000;
filter5[5][689] = 35'b00000010110011111101111101101000000;
filter5[5][690] = 35'b11111110111110111010100110011000000;
filter5[5][691] = 35'b00000000100011111111111100110101000;
filter5[5][692] = 35'b11111101101010101000110000111100000;
filter5[5][693] = 35'b00000000100000000100001011110010000;
filter5[5][694] = 35'b00000000001010001110010111011101100;
filter5[5][695] = 35'b00000101000000011100010000011000000;
filter5[5][696] = 35'b00000001101111000110011001100110000;
filter5[5][697] = 35'b00000000111000001110000100100000000;
filter5[5][698] = 35'b11111011110111010011100101101000000;
filter5[5][699] = 35'b00000001010101000101000101010010000;
filter5[5][700] = 35'b00000001111011100011011111101010000;
filter5[5][701] = 35'b00000101011010010101000000100000000;
filter5[5][702] = 35'b11111101110011100111001011101000000;
filter5[5][703] = 35'b00000011001000011001011111110000000;
filter5[5][704] = 35'b00000001110100100010100110110110000;
filter5[5][705] = 35'b11111111001000010101110111101111000;
filter5[5][706] = 35'b11111111100100101100001110110110100;
filter5[5][707] = 35'b11111100100101000010111000101000000;
filter5[5][708] = 35'b00000000011101011101111111110100000;
filter5[5][709] = 35'b00000000011000001110111001001110000;
filter5[5][710] = 35'b00000001010000101101010011011000000;
filter5[5][711] = 35'b11111111010001011101110110010001000;
filter5[5][712] = 35'b11111110001011001001011000110000000;
filter5[5][713] = 35'b11111110111111110110101001000000000;
filter5[5][714] = 35'b11111101110001101101100001001000000;
filter5[5][715] = 35'b11111101100010111001101101110100000;
filter5[5][716] = 35'b11111110011011011010001001000010000;
filter5[5][717] = 35'b00000001000000011101010011010010000;
filter5[5][718] = 35'b00000000111001010010001100101011000;
filter5[5][719] = 35'b11111110000101101100011101100000000;
filter5[5][720] = 35'b00000000000111000001101010110000110;
filter5[5][721] = 35'b00000000011001011010011111011101100;
filter5[5][722] = 35'b11111100101111110010001100111100000;
filter5[5][723] = 35'b00000010010011101001110010100000000;
filter5[5][724] = 35'b11111111011110111001110010101101000;
filter5[5][725] = 35'b00000010110000101010110011001100000;
filter5[5][726] = 35'b00000000100100111000101111100001000;
filter5[5][727] = 35'b11111100011110000000000111001000000;
filter5[5][728] = 35'b11111110101111111011011111010110000;
filter5[5][729] = 35'b11111110010001110100101101010110000;
filter5[5][730] = 35'b00000000011110110101011001101011000;
filter5[5][731] = 35'b00000001000010000000010110100000000;
filter5[5][732] = 35'b00000011000001001011111010111000000;
filter5[5][733] = 35'b00000000011001011100100011001011100;
filter5[5][734] = 35'b00000001110000001100100001011110000;
filter5[5][735] = 35'b11111100100110100100100000010100000;
filter5[5][736] = 35'b00000000001001001001111010010011100;
filter5[5][737] = 35'b11111110110100001110000010000100000;
filter5[5][738] = 35'b11111111010101001001110011001101000;
filter5[5][739] = 35'b11111110001111000100000001110010000;
filter5[5][740] = 35'b11111111100101111101101011011101100;
filter5[5][741] = 35'b11111111011101100100010000101001000;
filter5[5][742] = 35'b11111110101011010011110111001000000;
filter5[5][743] = 35'b00000000100111111110010001011110000;
filter5[5][744] = 35'b11111010011101001100000110011000000;
filter5[5][745] = 35'b00000001100101101000110110100010000;
filter5[5][746] = 35'b00000000001100010110101110111101110;
filter5[5][747] = 35'b00000000010110011001111111111111100;
filter5[5][748] = 35'b00000000010011110111101001000101100;
filter5[5][749] = 35'b00000010000111000110001000001100000;
filter5[5][750] = 35'b11111101101001100011001100111100000;
filter5[5][751] = 35'b00000011010110111100111110001000000;
filter5[5][752] = 35'b11111100111101000110101110111100000;
filter5[5][753] = 35'b11111100101110110110001100010100000;
filter5[5][754] = 35'b11111100101101000011010011110100000;
filter5[5][755] = 35'b11111110011001100001011010111100000;
filter5[5][756] = 35'b11111110000110100110010011011100000;
filter5[5][757] = 35'b00000011011001100001010000101000000;
filter5[5][758] = 35'b00000000100101011010001010000001000;
filter5[5][759] = 35'b00000100111001100010010011000000000;
filter5[5][760] = 35'b11111110000100000111110110100000000;
filter5[5][761] = 35'b11111100001000001011110000101000000;
filter5[5][762] = 35'b00000101001001001011111000011000000;
filter5[5][763] = 35'b11111111100110001100100000001101000;
filter5[5][764] = 35'b11111110000000101010111011110100000;
filter5[5][765] = 35'b00000001111000111010100111100100000;
filter5[5][766] = 35'b11111101100011100110100001110000000;
filter5[5][767] = 35'b00000000010010111111000000100101100;
filter5[5][768] = 35'b00000001101010011100001000000000000;
filter5[5][769] = 35'b00000010101000100000010100101000000;
filter5[5][770] = 35'b00000000010100000010110011000000100;
filter5[5][771] = 35'b00000011011001000010101001111100000;
filter5[5][772] = 35'b00000011001100111010010100100000000;
filter5[5][773] = 35'b00000001001011110000100110111010000;
filter5[5][774] = 35'b11111110010100111110101000011100000;
filter5[5][775] = 35'b11111011111011011001001101100000000;
filter5[5][776] = 35'b11111111000011101010011000001010000;
filter5[5][777] = 35'b11111110111101111110000101000010000;
filter5[5][778] = 35'b00000010010111111000111100010000000;
filter5[5][779] = 35'b00000000000100011000010010110110100;
filter5[5][780] = 35'b00000000101110011011011001100010000;
filter5[5][781] = 35'b00001000010100001011010111100000000;
filter5[5][782] = 35'b11111100001010001000110111010100000;
filter5[5][783] = 35'b00000000001101000011110111101011100;
filter5[5][784] = 35'b00000010000100010010101101110000000;
filter5[5][785] = 35'b11111111101110001111001100001011100;
filter5[5][786] = 35'b00000011001101100101111011011100000;
filter5[5][787] = 35'b00000001101001110000100111011010000;
filter5[5][788] = 35'b00000000110010100100110001010000000;
filter5[5][789] = 35'b11111101110000111110110011010000000;
filter5[5][790] = 35'b11111010110000001111101101000000000;
filter5[5][791] = 35'b00000000111010100100100101111000000;
filter5[5][792] = 35'b11111101110100101111100001111100000;
filter5[5][793] = 35'b00000001000011101010100101100100000;
filter5[5][794] = 35'b00000101000000101100010011101000000;
filter5[5][795] = 35'b11111111000111000011111101111100000;
filter5[5][796] = 35'b00000010011011011101100000010100000;
filter5[5][797] = 35'b11111100010000101010011001010100000;
filter5[5][798] = 35'b11111100011110100100010111010000000;
filter5[5][799] = 35'b11111100011101000001101010010000000;
filter5[5][800] = 35'b00000010111111011001100101111100000;
filter5[5][801] = 35'b11111111001000101110111111100100000;
filter5[5][802] = 35'b11111110001101101100001001100010000;
filter5[5][803] = 35'b00000001001010010101010111100110000;
filter5[5][804] = 35'b00000000101110011101010000011000000;
filter5[5][805] = 35'b11101110110001001111001110000000000;
filter5[5][806] = 35'b11111101000101111111110110111100000;
filter5[5][807] = 35'b11111001101110101101010101011000000;
filter5[5][808] = 35'b11111111110000000111111101110110110;
filter5[5][809] = 35'b11111110100110011000011110001110000;
filter5[5][810] = 35'b00000001100111100100111001011010000;
filter5[5][811] = 35'b11111100000110111001101100000000000;
filter5[5][812] = 35'b11110111111011011111111001110000000;
filter5[5][813] = 35'b11111011101001001000101001001000000;
filter5[5][814] = 35'b11111100011000000000001101011000000;
filter5[5][815] = 35'b00000010011001010001000100010000000;
filter5[5][816] = 35'b00000001111011101000110001100000000;
filter5[5][817] = 35'b00000001100110100100010010100110000;
filter5[5][818] = 35'b00000001100111011010001000100100000;
filter5[5][819] = 35'b00000000110110111000100111110000000;
filter5[5][820] = 35'b11111011110110101111011000001000000;
filter5[5][821] = 35'b00000000101011100011110100111111000;
filter5[5][822] = 35'b00000010100000101100111000100000000;
filter5[5][823] = 35'b00000001110111111011011101110010000;
filter5[5][824] = 35'b00000000000011110110000011011000111;
filter5[5][825] = 35'b00000000101000000001011100110100000;
filter5[5][826] = 35'b00000001111001011100011100110000000;
filter5[5][827] = 35'b11111101111100110101011010000000000;
filter5[5][828] = 35'b00000001101101000000111010110110000;
filter5[5][829] = 35'b11111111101010111100011011100101000;
filter5[5][830] = 35'b00000001000000100101010001100010000;
filter5[5][831] = 35'b00000010011111110101101001110100000;
filter5[5][832] = 35'b11111110001100000001101010000100000;
filter5[5][833] = 35'b11111100111111001111001001011000000;
filter5[5][834] = 35'b11111110101110000100111010100100000;
filter5[5][835] = 35'b11111110111010011010110100101010000;
filter5[5][836] = 35'b11111101110100111101101000001100000;
filter5[5][837] = 35'b11111111010001010000011010101000000;
filter5[5][838] = 35'b00000000000000000011101011100110011;
filter5[5][839] = 35'b11111111011001111111011110110100000;
filter5[5][840] = 35'b00000000011000000101101000110001000;
filter5[5][841] = 35'b11111101011000101001010110111000000;
filter5[5][842] = 35'b11111100110001000001010110010100000;
filter5[5][843] = 35'b11111110111100111000111100001100000;
filter5[5][844] = 35'b00000001100110010100111010000100000;
filter5[5][845] = 35'b00000000011101011110101110000101100;
filter5[5][846] = 35'b11111110110010101110001000100000000;
filter5[5][847] = 35'b11111111100110100101001011010110100;
filter5[5][848] = 35'b11111111011111101010011000011011000;
filter5[5][849] = 35'b11111101001110101010010001001100000;
filter5[5][850] = 35'b11111101110110101110110111100100000;
filter5[5][851] = 35'b11111111111100110000010001111011011;
filter5[5][852] = 35'b00000000011001010101110011100001000;
filter5[5][853] = 35'b00000110111100110111101101101000000;
filter5[5][854] = 35'b00000001100001100111101001011010000;
filter5[5][855] = 35'b11111010110100110001111111101000000;
filter5[5][856] = 35'b11111101011111100111110000110000000;
filter5[5][857] = 35'b11111101000100101110100101110000000;
filter5[5][858] = 35'b11111111000010110010011100111101000;
filter5[5][859] = 35'b11111111011001010101101111011011000;
filter5[5][860] = 35'b00000100000000101101111111010000000;
filter5[5][861] = 35'b11111110011110100101010111000010000;
filter5[5][862] = 35'b11111110111100110011101001110010000;
filter5[5][863] = 35'b11111010100110010000110110011000000;
filter5[5][864] = 35'b11111101000111100100100011100100000;
filter5[5][865] = 35'b11111110111101000010011101100110000;
filter5[5][866] = 35'b00000001111011001101011111001010000;
filter5[5][867] = 35'b11111110010101111011010100111000000;
filter5[5][868] = 35'b11111111110010100000101110101111100;
filter5[5][869] = 35'b00000000111111110010100011000100000;
filter5[5][870] = 35'b00000001111010001111000000101100000;
filter5[5][871] = 35'b00000010111001001011101111110100000;
filter5[5][872] = 35'b11111101000111100000100110001000000;
filter5[5][873] = 35'b00000001010010010101010011001100000;
filter5[5][874] = 35'b00000010010000111101000001010000000;
filter5[5][875] = 35'b00000001100110000110000010100110000;
filter5[5][876] = 35'b00000001001110000011110001000010000;
filter5[5][877] = 35'b00000001010011100101110011111000000;
filter5[5][878] = 35'b11111111011000001000000111111000000;
filter5[5][879] = 35'b11111011000011111011101110100000000;
filter5[5][880] = 35'b11111101000000010011100101011100000;
filter5[5][881] = 35'b00000001101010011001110111000100000;
filter5[5][882] = 35'b11111001110101001000110111001000000;
filter5[5][883] = 35'b00000000000110101111011101111110111;
filter5[5][884] = 35'b00000001101110110110011001000100000;
filter5[5][885] = 35'b00000011011101111111000001101000000;
filter5[5][886] = 35'b00000000111111010010111001101110000;
filter5[5][887] = 35'b00000011011000110101111010000000000;
filter5[5][888] = 35'b11111101000000100110010011111100000;
filter5[5][889] = 35'b11111001110101101001100101100000000;
filter5[5][890] = 35'b11111101010100001110100111001100000;
filter5[5][891] = 35'b11111100001001101001100010001000000;
filter5[5][892] = 35'b00000001011000111010001001011010000;
filter5[5][893] = 35'b11111111001111101000110010100011000;
filter5[5][894] = 35'b11111111000110011111001000001010000;
filter5[5][895] = 35'b00000001011010000000100101000100000;
filter5[5][896] = 35'b00000011011010001000110111110000000;
filter5[5][897] = 35'b00000001010010000111011101100100000;
filter5[5][898] = 35'b11111011111001111111010010101000000;
filter5[5][899] = 35'b11110000111111000000110110000000000;
filter5[5][900] = 35'b00000101100100010110110110110000000;
filter5[5][901] = 35'b00000011101011000101001011100100000;
filter5[5][902] = 35'b00000101100000101000100111101000000;
filter5[5][903] = 35'b00000010110100111111000110101000000;
filter5[5][904] = 35'b00001000010000101000100101010000000;
filter5[5][905] = 35'b11111100100000101110111110001100000;
filter5[5][906] = 35'b11111000001100011011101010110000000;
filter5[5][907] = 35'b11111111101101011001100110011100100;
filter5[5][908] = 35'b11111111011100100001100010110100000;
filter5[5][909] = 35'b00000100110000010011001001011000000;
filter5[5][910] = 35'b00000100100000010111000101100000000;
filter5[5][911] = 35'b11111110100111111010100101001100000;
filter5[5][912] = 35'b11111001110010001000010101111000000;
filter5[5][913] = 35'b11110110111111101010111110000000000;
filter5[5][914] = 35'b00000000101101011110101011000011000;
filter5[5][915] = 35'b11111110010000100101110010100110000;
filter5[5][916] = 35'b00000001000000101110100100000110000;
filter5[5][917] = 35'b00000001101100100000001001101110000;
filter5[5][918] = 35'b11111110111101110110010010010100000;
filter5[5][919] = 35'b11110101110000111011101000000000000;
filter5[5][920] = 35'b00000010011000001000000000110100000;
filter5[5][921] = 35'b11111111000100001110100001111000000;
filter5[5][922] = 35'b00000011100111100101110110100000000;
filter5[5][923] = 35'b11111111111110000111100100110101100;
filter5[5][924] = 35'b00000001101001100111101100010100000;
filter5[5][925] = 35'b00000010100111110100110001110000000;
filter5[5][926] = 35'b11111111000011110111001000111101000;
filter5[5][927] = 35'b11111110111001000000100111101100000;
filter5[5][928] = 35'b11111100000100100110001111011100000;
filter5[5][929] = 35'b11111111101110101010110111011011000;
filter5[5][930] = 35'b00000001100111101100000111101010000;
filter5[5][931] = 35'b11111111000001001110111111010100000;
filter5[5][932] = 35'b11111111000011110000000001110010000;
filter5[5][933] = 35'b11111111100010001011111000011101000;
filter5[5][934] = 35'b11111100100011101101010010111100000;
filter5[5][935] = 35'b00000110000111011011001011010000000;
filter5[5][936] = 35'b11111101010111001111101100001100000;
filter5[5][937] = 35'b11111101100100110110011100111100000;
filter5[5][938] = 35'b11111110001010110010101000111010000;
filter5[5][939] = 35'b11111111010001011000110100010011000;
filter5[5][940] = 35'b00000000100111101000001001110010000;
filter5[5][941] = 35'b00000010001100111110101111100000000;
filter5[5][942] = 35'b00000001110100011110100101100010000;
filter5[5][943] = 35'b00000100011100001001011011111000000;
filter5[5][944] = 35'b11111011011111010111110011011000000;
filter5[5][945] = 35'b11111010101001111011101100001000000;
filter5[5][946] = 35'b11111100111001110110000010101100000;
filter5[5][947] = 35'b11111101100010100001000100110000000;
filter5[5][948] = 35'b00000100010001001111111100111000000;
filter5[5][949] = 35'b00000001000011111100101011001000000;
filter5[5][950] = 35'b11111110110111101000100110010000000;
filter5[5][951] = 35'b00000111111011111111000011100000000;
filter5[5][952] = 35'b11111011011110101110101000010000000;
filter5[5][953] = 35'b11110101000101000100000010110000000;
filter5[5][954] = 35'b00000111000111011001011100100000000;
filter5[5][955] = 35'b11111100000101001001110100110000000;
filter5[5][956] = 35'b11111101000111110101000000100000000;
filter5[5][957] = 35'b11111101010101101111111110111000000;
filter5[5][958] = 35'b11111011111111100001110001011000000;
filter5[5][959] = 35'b00000111011000000001001100000000000;
filter5[5][960] = 35'b11111101101011000111100001001100000;
filter5[5][961] = 35'b00000100111001101010000100010000000;
filter5[5][962] = 35'b11111001000001001001101111010000000;
filter5[5][963] = 35'b11110101000100101110010000010000000;
filter5[5][964] = 35'b00000001011111110111110100100010000;
filter5[5][965] = 35'b00000100100010000100011111100000000;
filter5[5][966] = 35'b00000011111010010001001111010100000;
filter5[5][967] = 35'b00000111000010011010001110011000000;
filter5[5][968] = 35'b11111101111001101101001010001000000;
filter5[5][969] = 35'b11111000111111000011111110001000000;
filter5[5][970] = 35'b11110011111011111000111111000000000;
filter5[5][971] = 35'b11111101100100011010100100011000000;
filter5[5][972] = 35'b00000001111111010001001010110000000;
filter5[5][973] = 35'b00000010100101101001000111100000000;
filter5[5][974] = 35'b00000010101100010010001100111000000;
filter5[5][975] = 35'b00000000110010000111000111110110000;
filter5[5][976] = 35'b11110101000011100000001000100000000;
filter5[5][977] = 35'b11111100100001101001110111101100000;
filter5[5][978] = 35'b11111110110100000110100101111010000;
filter5[5][979] = 35'b00000000100010011001000100010001000;
filter5[5][980] = 35'b11111111011111110001111001110011000;
filter5[5][981] = 35'b00000000000001000101100100110001011;
filter5[5][982] = 35'b11111111100001001011010111010010100;
filter5[5][983] = 35'b00000000101011111010000011110100000;
filter5[5][984] = 35'b11110001101111000101100110000000000;
filter5[5][985] = 35'b11111011010010000011011101001000000;
filter5[5][986] = 35'b00000011000011001000111111101000000;
filter5[5][987] = 35'b00000011110101000011111010101000000;
filter5[5][988] = 35'b11111101011101100100011100011000000;
filter5[5][989] = 35'b11111111010010011100011000000001000;
filter5[5][990] = 35'b11111110011010000111011011100100000;
filter5[5][991] = 35'b00000110001111011100110000110000000;
filter5[5][992] = 35'b11110101001100110011100100100000000;
filter5[5][993] = 35'b11110111111001010001111101010000000;
filter5[5][994] = 35'b11110111011000011001011110000000000;
filter5[5][995] = 35'b11111110101000000000111011111110000;
filter5[5][996] = 35'b00000000101100101011111000000011000;
filter5[5][997] = 35'b00000001101100011101100100001000000;
filter5[5][998] = 35'b00000100010000001010101101001000000;
filter5[5][999] = 35'b11111100011100000010000110011100000;
filter5[5][1000] = 35'b11111100001100001100010001101000000;
filter5[5][1001] = 35'b00000110011011110010110000010000000;
filter5[5][1002] = 35'b11110011100011110100101111110000000;
filter5[5][1003] = 35'b11111101011010000110001110101100000;
filter5[5][1004] = 35'b00000001111110101110101110000110000;
filter5[5][1005] = 35'b00000010100000000111111001101100000;
filter5[5][1006] = 35'b00000101001100111111100101000000000;
filter5[5][1007] = 35'b11111100001111101011111001001000000;
filter5[5][1008] = 35'b11111010010001010000000011101000000;
filter5[5][1009] = 35'b11110010010110111001000100010000000;
filter5[5][1010] = 35'b11110110001000101101000111100000000;
filter5[5][1011] = 35'b11111011100110100101110011111000000;
filter5[5][1012] = 35'b00000000001010011101100011001110100;
filter5[5][1013] = 35'b00000010000100011000010110110100000;
filter5[5][1014] = 35'b00000010001011001000101000010000000;
filter5[5][1015] = 35'b11111111111000010101110101110100001;
filter5[5][1016] = 35'b11111111110100000000001111010100000;
filter5[5][1017] = 35'b11111110010001010110100010001100000;
filter5[5][1018] = 35'b11111000011110010010100101111000000;
filter5[5][1019] = 35'b00000000100000101111001110100000000;
filter5[5][1020] = 35'b00000000010001011110111101010111000;
filter5[5][1021] = 35'b11111010010100010000011011110000000;
filter5[5][1022] = 35'b00000001111010111000000010111010000;
filter5[5][1023] = 35'b00000111000101000011101101010000000;
filter5[6][0] = 35'b00000010000101011001010010001000000;
filter5[6][1] = 35'b00000110111111011111111010000000000;
filter5[6][2] = 35'b00000011011000111000000110111100000;
filter5[6][3] = 35'b11111001111001101110111000001000000;
filter5[6][4] = 35'b00000000111010011101000111010000000;
filter5[6][5] = 35'b11111110011000010011110101000110000;
filter5[6][6] = 35'b11111101110111110011011011111000000;
filter5[6][7] = 35'b11110111000000010101000101100000000;
filter5[6][8] = 35'b00000010011001000000100010110000000;
filter5[6][9] = 35'b11111101101001001001011001000000000;
filter5[6][10] = 35'b00000010110010110001110000111100000;
filter5[6][11] = 35'b00000110111011010111110100110000000;
filter5[6][12] = 35'b11111111110111011000110110110010010;
filter5[6][13] = 35'b11111111100100110101110001100001000;
filter5[6][14] = 35'b00000101001110110100110011100000000;
filter5[6][15] = 35'b11110111011100011001000000000000000;
filter5[6][16] = 35'b00000010010101000001011000011100000;
filter5[6][17] = 35'b11111111111110110100101100001000100;
filter5[6][18] = 35'b00000110000010101001000111000000000;
filter5[6][19] = 35'b11111110111001101110110010000110000;
filter5[6][20] = 35'b11111110101000100011100110110110000;
filter5[6][21] = 35'b00000001000011000010111001001110000;
filter5[6][22] = 35'b11111111111110010101010011001011010;
filter5[6][23] = 35'b11111011100001001001011110001000000;
filter5[6][24] = 35'b11111101000111110001011001010100000;
filter5[6][25] = 35'b11111101100111101110101011111100000;
filter5[6][26] = 35'b00000010000111010100001100101100000;
filter5[6][27] = 35'b00000000010011011110101001100111000;
filter5[6][28] = 35'b11111110011011010011001011011110000;
filter5[6][29] = 35'b00000000011101011010010000011100000;
filter5[6][30] = 35'b00001000111110111001010011100000000;
filter5[6][31] = 35'b00000011001011001110100001100100000;
filter5[6][32] = 35'b11111011100111101111001100001000000;
filter5[6][33] = 35'b11111101110000111010110000011000000;
filter5[6][34] = 35'b11111110000000110001111110010110000;
filter5[6][35] = 35'b11111101011110011101110100000100000;
filter5[6][36] = 35'b11111110100010010010101000010000000;
filter5[6][37] = 35'b11111101101010100001100011110000000;
filter5[6][38] = 35'b00000000100001001100000101111111000;
filter5[6][39] = 35'b00000110110000000111011101111000000;
filter5[6][40] = 35'b11111100101011001110010100001000000;
filter5[6][41] = 35'b00000001100001001010000010000010000;
filter5[6][42] = 35'b11111110100110100001001101010100000;
filter5[6][43] = 35'b00000000101000100100010010100011000;
filter5[6][44] = 35'b00000101010010010111011100011000000;
filter5[6][45] = 35'b00000010010010001000111001111100000;
filter5[6][46] = 35'b11111101111000100100100011001000000;
filter5[6][47] = 35'b11111110001010000100000011001010000;
filter5[6][48] = 35'b11111001110110000011011000010000000;
filter5[6][49] = 35'b00000001111101111101010111000000000;
filter5[6][50] = 35'b00000000011010000011010010011110100;
filter5[6][51] = 35'b00000001100010001100001111010000000;
filter5[6][52] = 35'b00001001000111001100101001000000000;
filter5[6][53] = 35'b11111001100000001010011100001000000;
filter5[6][54] = 35'b11111100111110101000111111111100000;
filter5[6][55] = 35'b00000001110110110101000111101010000;
filter5[6][56] = 35'b00000100101101011100000010110000000;
filter5[6][57] = 35'b11110111111101010100111111100000000;
filter5[6][58] = 35'b00000010110011000110101100011000000;
filter5[6][59] = 35'b00000011101111011000010100101100000;
filter5[6][60] = 35'b11111100011100100111001100000100000;
filter5[6][61] = 35'b11111111000101111011000001011001000;
filter5[6][62] = 35'b11111011000000100011010111100000000;
filter5[6][63] = 35'b11111001010000101011000001001000000;
filter5[6][64] = 35'b11111111011110111111010011000101000;
filter5[6][65] = 35'b00000010101001010001111001000100000;
filter5[6][66] = 35'b11111111111001101100101000011101100;
filter5[6][67] = 35'b11111010011010110000010100110000000;
filter5[6][68] = 35'b11111100000000110110101101011100000;
filter5[6][69] = 35'b00000010101010000001010101100100000;
filter5[6][70] = 35'b00000001100110011110111111100000000;
filter5[6][71] = 35'b11111000010011001111000111100000000;
filter5[6][72] = 35'b00000010001010110011001110100100000;
filter5[6][73] = 35'b11111001110100001110011101011000000;
filter5[6][74] = 35'b11111010000010110110101111110000000;
filter5[6][75] = 35'b00000001101101011010001110001100000;
filter5[6][76] = 35'b11111101011100010011001011011000000;
filter5[6][77] = 35'b00000001001110110101010100010100000;
filter5[6][78] = 35'b11111110101100100011100110000010000;
filter5[6][79] = 35'b11111101110111101011010111010100000;
filter5[6][80] = 35'b00000100101010011010101101010000000;
filter5[6][81] = 35'b11111111011111111011101110001111000;
filter5[6][82] = 35'b00000010000001101111010101011100000;
filter5[6][83] = 35'b11111011110010010010100110010000000;
filter5[6][84] = 35'b11111111101100010101000101101100100;
filter5[6][85] = 35'b00000000111010111010110100100000000;
filter5[6][86] = 35'b11111111001000100110111000011110000;
filter5[6][87] = 35'b11111111000011101111000110111111000;
filter5[6][88] = 35'b11111110000010000010100010111010000;
filter5[6][89] = 35'b00000000001001100000000100100010100;
filter5[6][90] = 35'b00000011100100001110000011110100000;
filter5[6][91] = 35'b00000010011011010100000110001000000;
filter5[6][92] = 35'b00000001100100100101111000111110000;
filter5[6][93] = 35'b00000011100011110001101001011000000;
filter5[6][94] = 35'b11111111101101111101101111011111100;
filter5[6][95] = 35'b00000000001110011111011010000001110;
filter5[6][96] = 35'b11111011101011011001101010101000000;
filter5[6][97] = 35'b11111110111000011100101101100100000;
filter5[6][98] = 35'b00000010010101011001001110010000000;
filter5[6][99] = 35'b11111101110000011101111110000100000;
filter5[6][100] = 35'b00000000000101011101000111001111101;
filter5[6][101] = 35'b11111111001001101110011100100010000;
filter5[6][102] = 35'b11111111100001011001111100101111100;
filter5[6][103] = 35'b11111110100101000100011000100110000;
filter5[6][104] = 35'b11111101101100011010101001000100000;
filter5[6][105] = 35'b11111101001010001000100110101000000;
filter5[6][106] = 35'b11111111100011011001010101110100000;
filter5[6][107] = 35'b00000000001100101101111111001100100;
filter5[6][108] = 35'b00000000011001001110011000110001100;
filter5[6][109] = 35'b11111110101011001011001110100000000;
filter5[6][110] = 35'b00000010111010111110100001001000000;
filter5[6][111] = 35'b11111110010011000111001010010100000;
filter5[6][112] = 35'b00000000011101011100101110101101000;
filter5[6][113] = 35'b11111101010110010111000001111000000;
filter5[6][114] = 35'b11111101100110001101011111010100000;
filter5[6][115] = 35'b00000010001100000111011101110100000;
filter5[6][116] = 35'b00000000110111010000110110100000000;
filter5[6][117] = 35'b11111111100110010011011101001110100;
filter5[6][118] = 35'b00000011111110011001000110000000000;
filter5[6][119] = 35'b00000010100011010111100100010100000;
filter5[6][120] = 35'b00000101011001110111001011010000000;
filter5[6][121] = 35'b11110001111111100000101000110000000;
filter5[6][122] = 35'b00000010111000000001000001100000000;
filter5[6][123] = 35'b00000000010011010001100111110001000;
filter5[6][124] = 35'b00000010110101010111010010101100000;
filter5[6][125] = 35'b11111110010000110010101010010110000;
filter5[6][126] = 35'b00001001011100011111111110000000000;
filter5[6][127] = 35'b00000001101101000111001011101000000;
filter5[6][128] = 35'b11111110000010111010111001000100000;
filter5[6][129] = 35'b11111111111011110100110110010101011;
filter5[6][130] = 35'b11111000100000001010000101000000000;
filter5[6][131] = 35'b11101001101000110110111000100000000;
filter5[6][132] = 35'b11111010110001100011011010000000000;
filter5[6][133] = 35'b00000101110010101101001100000000000;
filter5[6][134] = 35'b00001000100011001000000100010000000;
filter5[6][135] = 35'b11111001010010001111000100111000000;
filter5[6][136] = 35'b11111011001111011011001000110000000;
filter5[6][137] = 35'b11101110001011010010100111100000000;
filter5[6][138] = 35'b11110111010010011000110110000000000;
filter5[6][139] = 35'b00000100011101111000101100101000000;
filter5[6][140] = 35'b11111110110111010100110110111100000;
filter5[6][141] = 35'b00000000011101010110010111101001100;
filter5[6][142] = 35'b11111110101000101101010010110010000;
filter5[6][143] = 35'b11111111110111000111010110011011000;
filter5[6][144] = 35'b00000000111010111010000111000011000;
filter5[6][145] = 35'b11111000100110101011110100011000000;
filter5[6][146] = 35'b00000101110011001111001110011000000;
filter5[6][147] = 35'b00000001011010001100110011000110000;
filter5[6][148] = 35'b00000010001101011001000010000100000;
filter5[6][149] = 35'b11111110011001010110111101101010000;
filter5[6][150] = 35'b11111111101101000010110110111111000;
filter5[6][151] = 35'b00000001001011101111000101011000000;
filter5[6][152] = 35'b11111101011000100110111001111000000;
filter5[6][153] = 35'b00000000100000011010100010111000000;
filter5[6][154] = 35'b00000100110111111100011100001000000;
filter5[6][155] = 35'b00000011001111001000100110111100000;
filter5[6][156] = 35'b00000100110011011011001110101000000;
filter5[6][157] = 35'b11111111000101101110001000011100000;
filter5[6][158] = 35'b11111101101010100110010110010000000;
filter5[6][159] = 35'b11111101011111101010011010011100000;
filter5[6][160] = 35'b00000010011110101010100001010000000;
filter5[6][161] = 35'b11110110111001011110011000110000000;
filter5[6][162] = 35'b11111001001000111010000100110000000;
filter5[6][163] = 35'b11111010011010001111010001011000000;
filter5[6][164] = 35'b11111100110101111011010010001100000;
filter5[6][165] = 35'b00000001011010111010111100100000000;
filter5[6][166] = 35'b00000000010110001110101110000111100;
filter5[6][167] = 35'b11110110011000111101100110000000000;
filter5[6][168] = 35'b11110101000101001100000010100000000;
filter5[6][169] = 35'b11111011100101010011111111110000000;
filter5[6][170] = 35'b11111101100101100110101011000000000;
filter5[6][171] = 35'b11111010000110000000110100101000000;
filter5[6][172] = 35'b11111000010010001101001000001000000;
filter5[6][173] = 35'b00000001110001100011110111010110000;
filter5[6][174] = 35'b11111110111001111111010111001000000;
filter5[6][175] = 35'b11110110011100100110101010000000000;
filter5[6][176] = 35'b11110111101001010011011010100000000;
filter5[6][177] = 35'b11110101011111111100011011100000000;
filter5[6][178] = 35'b11111010011000010100110100111000000;
filter5[6][179] = 35'b11110100101101111001101011100000000;
filter5[6][180] = 35'b11101011001100100101111101100000000;
filter5[6][181] = 35'b00000110011100100011110011100000000;
filter5[6][182] = 35'b00010010000010000000101001100000000;
filter5[6][183] = 35'b11101011101101111100100001000000000;
filter5[6][184] = 35'b00000111100000110111111001110000000;
filter5[6][185] = 35'b11111110011011110011100100001000000;
filter5[6][186] = 35'b00000011110000001100101110100000000;
filter5[6][187] = 35'b11111011111110011011100110011000000;
filter5[6][188] = 35'b00000001000001101111001011110110000;
filter5[6][189] = 35'b11110111000010101001000010110000000;
filter5[6][190] = 35'b11111111101101101111001010011001100;
filter5[6][191] = 35'b11100100100011111001001110000000000;
filter5[6][192] = 35'b11111111100101000010111111000011000;
filter5[6][193] = 35'b00000000001011100011011101110101100;
filter5[6][194] = 35'b11111011110110000111010101110000000;
filter5[6][195] = 35'b11110110101100000111010100110000000;
filter5[6][196] = 35'b11111001100111111000111010110000000;
filter5[6][197] = 35'b11110100110101111101001110000000000;
filter5[6][198] = 35'b11110110101110000100101101110000000;
filter5[6][199] = 35'b11101100111000010011001010000000000;
filter5[6][200] = 35'b11110110001001111101010110110000000;
filter5[6][201] = 35'b00000110000110000010101001101000000;
filter5[6][202] = 35'b11110000001000001011010111100000000;
filter5[6][203] = 35'b11111000001110100001110001010000000;
filter5[6][204] = 35'b00000001111110010000101011100010000;
filter5[6][205] = 35'b00000110011111001011111010011000000;
filter5[6][206] = 35'b11111101011000111011111001100100000;
filter5[6][207] = 35'b00001001000110010010010001110000000;
filter5[6][208] = 35'b11111111101001010101111011001110100;
filter5[6][209] = 35'b00000000010010101101000110110101100;
filter5[6][210] = 35'b11111010101101000010111110101000000;
filter5[6][211] = 35'b11111001111100111111101000100000000;
filter5[6][212] = 35'b00000000110110101110101011010111000;
filter5[6][213] = 35'b00000001010110000110101001101000000;
filter5[6][214] = 35'b00000010111010001110011010110000000;
filter5[6][215] = 35'b00000010001011000101001001010000000;
filter5[6][216] = 35'b11111011111110011111101100110000000;
filter5[6][217] = 35'b11110001111111000010000001110000000;
filter5[6][218] = 35'b11111110110111010110000100000110000;
filter5[6][219] = 35'b00000011111110010100001011111000000;
filter5[6][220] = 35'b00000000011111111010100010001001000;
filter5[6][221] = 35'b00000001000000101001100111111100000;
filter5[6][222] = 35'b11111111101001001011000101000101000;
filter5[6][223] = 35'b11111100100011011101111101001000000;
filter5[6][224] = 35'b11111100100001011110000001111000000;
filter5[6][225] = 35'b11111000111000001100011011110000000;
filter5[6][226] = 35'b11111111110000101001110111101011110;
filter5[6][227] = 35'b11111110000110000111110010101110000;
filter5[6][228] = 35'b11111111000001111011010100101011000;
filter5[6][229] = 35'b00000001011100001111111111110010000;
filter5[6][230] = 35'b11111111101010010000100010110100000;
filter5[6][231] = 35'b00000010110010010101110111100000000;
filter5[6][232] = 35'b11101001000110111011100101000000000;
filter5[6][233] = 35'b00000100101001111111100111110000000;
filter5[6][234] = 35'b11111011100111011011001101001000000;
filter5[6][235] = 35'b11111110011000110111010000100000000;
filter5[6][236] = 35'b11111111111000100110000101101001101;
filter5[6][237] = 35'b00000010111000010101000000100000000;
filter5[6][238] = 35'b11111101011001100000010000000100000;
filter5[6][239] = 35'b11111101101111110111111111001100000;
filter5[6][240] = 35'b11111101110011100010101100100000000;
filter5[6][241] = 35'b00000011011101000100001000101000000;
filter5[6][242] = 35'b11111011010111000011001110100000000;
filter5[6][243] = 35'b11111100000100011100100011001100000;
filter5[6][244] = 35'b00000001000110110100010001100000000;
filter5[6][245] = 35'b00000100010110000010010101011000000;
filter5[6][246] = 35'b11111110101011000100111010100010000;
filter5[6][247] = 35'b00000100011101111101011110100000000;
filter5[6][248] = 35'b11111000111111100111000100111000000;
filter5[6][249] = 35'b11111111101000110110000101111000000;
filter5[6][250] = 35'b11111001001001011101000100110000000;
filter5[6][251] = 35'b00000000111101000000100111000001000;
filter5[6][252] = 35'b11111110011000110000000011100100000;
filter5[6][253] = 35'b00000010110101111101110100100000000;
filter5[6][254] = 35'b00000010001010010100000111010100000;
filter5[6][255] = 35'b00000010010011101010100110100100000;
filter5[6][256] = 35'b00000100000001011100001000100000000;
filter5[6][257] = 35'b11111111111111000011010001101010001;
filter5[6][258] = 35'b11111111001001011000001010101010000;
filter5[6][259] = 35'b11110100110011001101001000010000000;
filter5[6][260] = 35'b11111011100111000111110000100000000;
filter5[6][261] = 35'b11110100101010111001010010110000000;
filter5[6][262] = 35'b11110110000101110101001010110000000;
filter5[6][263] = 35'b11111001110001101000110011111000000;
filter5[6][264] = 35'b11111011101111000011010111001000000;
filter5[6][265] = 35'b11111011110111001110101010110000000;
filter5[6][266] = 35'b11110010001100110110010100000000000;
filter5[6][267] = 35'b11111111011001010100000101111101000;
filter5[6][268] = 35'b00001010010000100110001110110000000;
filter5[6][269] = 35'b11111011110010001011010000100000000;
filter5[6][270] = 35'b00000100111001111000100111111000000;
filter5[6][271] = 35'b00000101001000101010100101000000000;
filter5[6][272] = 35'b00000100101011100101111101100000000;
filter5[6][273] = 35'b11110011010010111010110011110000000;
filter5[6][274] = 35'b11111010000001011101011100100000000;
filter5[6][275] = 35'b11111111000110000011000111000010000;
filter5[6][276] = 35'b00000100100011101101110000010000000;
filter5[6][277] = 35'b00000000011000010111100010011110100;
filter5[6][278] = 35'b00000001001101011101100110001100000;
filter5[6][279] = 35'b11111101000000011111110010001000000;
filter5[6][280] = 35'b11111001011011101011110101111000000;
filter5[6][281] = 35'b11110011110010010000110001000000000;
filter5[6][282] = 35'b11111100111101110011000001011100000;
filter5[6][283] = 35'b11111111111101110101010010111101110;
filter5[6][284] = 35'b11111101011010001000000000101100000;
filter5[6][285] = 35'b11111111110100111011101001011110100;
filter5[6][286] = 35'b11111101000000110101110100000100000;
filter5[6][287] = 35'b00000010000011111101011111001000000;
filter5[6][288] = 35'b11110111110011000010011110110000000;
filter5[6][289] = 35'b11111100011010101101111010100000000;
filter5[6][290] = 35'b11111101101001000011101100111100000;
filter5[6][291] = 35'b00000011000000101110110010001000000;
filter5[6][292] = 35'b11111101110101011100111001100100000;
filter5[6][293] = 35'b11111101101111001101100000110000000;
filter5[6][294] = 35'b11111111111011110001111101111100001;
filter5[6][295] = 35'b00000001111010011000101100110010000;
filter5[6][296] = 35'b00000010000010001110110000011000000;
filter5[6][297] = 35'b11111101100101000101111010010000000;
filter5[6][298] = 35'b11111011001001001010000000011000000;
filter5[6][299] = 35'b11111100100101100011011010010100000;
filter5[6][300] = 35'b00000010101100111000010111011000000;
filter5[6][301] = 35'b00000010111000111100010100011100000;
filter5[6][302] = 35'b00000010111111110110110011011000000;
filter5[6][303] = 35'b00000001000101001111110100001010000;
filter5[6][304] = 35'b00000100000001011000100110101000000;
filter5[6][305] = 35'b11111010111000111010001110111000000;
filter5[6][306] = 35'b11111101110111011111100111001000000;
filter5[6][307] = 35'b11111010010101111110011110010000000;
filter5[6][308] = 35'b00000011101111001011001110111000000;
filter5[6][309] = 35'b11111111000101001011001011010000000;
filter5[6][310] = 35'b11111110101001010111010100001010000;
filter5[6][311] = 35'b00000000010101010001100111001100100;
filter5[6][312] = 35'b11101001110010010101001010000000000;
filter5[6][313] = 35'b11110010000010101011010011010000000;
filter5[6][314] = 35'b00000101101111110001011111100000000;
filter5[6][315] = 35'b11111010101000101101111011010000000;
filter5[6][316] = 35'b00000010001110111011111011000000000;
filter5[6][317] = 35'b00000110010100100110011010001000000;
filter5[6][318] = 35'b11111111011000000011001111111011000;
filter5[6][319] = 35'b00000110101000010101001100100000000;
filter5[6][320] = 35'b11111011100110010000011110000000000;
filter5[6][321] = 35'b00000000000110000100000000010101001;
filter5[6][322] = 35'b11111111101011100010001000010010100;
filter5[6][323] = 35'b11110111000000011111010001100000000;
filter5[6][324] = 35'b00000010110010001010111110101000000;
filter5[6][325] = 35'b00001000110111110110000000010000000;
filter5[6][326] = 35'b11111111010101100101111100001001000;
filter5[6][327] = 35'b11110110011110010101110110000000000;
filter5[6][328] = 35'b11110111001110001100010101010000000;
filter5[6][329] = 35'b11111101101010101110101010010100000;
filter5[6][330] = 35'b11111011111100001001101001000000000;
filter5[6][331] = 35'b11111101001110110110100101101000000;
filter5[6][332] = 35'b00000000000110010001011111111011010;
filter5[6][333] = 35'b00000101100001010010000110100000000;
filter5[6][334] = 35'b00000000000001010101111010111101110;
filter5[6][335] = 35'b11111011110101111010110001011000000;
filter5[6][336] = 35'b11111111101110111111001010000111100;
filter5[6][337] = 35'b11111111011001001001111011000011000;
filter5[6][338] = 35'b00000010000111001000011011011100000;
filter5[6][339] = 35'b00000001000010010011100010111100000;
filter5[6][340] = 35'b11111110101001000110001111100100000;
filter5[6][341] = 35'b00000001110011011101100000110010000;
filter5[6][342] = 35'b11111111000001011110101110000000000;
filter5[6][343] = 35'b11111111111001110001001111011000011;
filter5[6][344] = 35'b00000000001011111101101011110111100;
filter5[6][345] = 35'b11111101111010011011010100110100000;
filter5[6][346] = 35'b00000000001001010101001011000010010;
filter5[6][347] = 35'b00000001111000101110110001001100000;
filter5[6][348] = 35'b11111110010111001111111011100000000;
filter5[6][349] = 35'b11111111100101101011011001010111100;
filter5[6][350] = 35'b11111111000001011110101111101100000;
filter5[6][351] = 35'b11111101111100101101111001101100000;
filter5[6][352] = 35'b11111111000110001010100000001001000;
filter5[6][353] = 35'b00000000010101101011010111000110000;
filter5[6][354] = 35'b00000000110000001110001101111011000;
filter5[6][355] = 35'b11111111001001110110101010101010000;
filter5[6][356] = 35'b11111110101010110010001111101100000;
filter5[6][357] = 35'b00000000111000101010110111001101000;
filter5[6][358] = 35'b11111111000101011111000110110000000;
filter5[6][359] = 35'b00000000111101010010011000000101000;
filter5[6][360] = 35'b11111011111100000100010000100000000;
filter5[6][361] = 35'b00000001101110100110100100111000000;
filter5[6][362] = 35'b11111101001101111111011010100000000;
filter5[6][363] = 35'b00000000111100010010011011000011000;
filter5[6][364] = 35'b00000010010111001011001100000000000;
filter5[6][365] = 35'b00000001100100011111110011010010000;
filter5[6][366] = 35'b00000001101000001011010110101000000;
filter5[6][367] = 35'b00000000001100001000101111101100010;
filter5[6][368] = 35'b11111011010101101101110000010000000;
filter5[6][369] = 35'b11111110110011110101101011111000000;
filter5[6][370] = 35'b00000001110110110110011011101010000;
filter5[6][371] = 35'b11111111100010000010100100110010100;
filter5[6][372] = 35'b00000000100001001100001000010111000;
filter5[6][373] = 35'b11111101001101101001111111000000000;
filter5[6][374] = 35'b00000010101011010010101000011100000;
filter5[6][375] = 35'b00000011011001101100011001101100000;
filter5[6][376] = 35'b00000111010010000100010110000000000;
filter5[6][377] = 35'b11111011000111000110110001010000000;
filter5[6][378] = 35'b11111111110001110101100001111101000;
filter5[6][379] = 35'b11111111001000010100100011011110000;
filter5[6][380] = 35'b00000001001001010001101000111010000;
filter5[6][381] = 35'b00000010110100101100101010010100000;
filter5[6][382] = 35'b00000011010100011100100011100000000;
filter5[6][383] = 35'b11111111111011111100111001101101100;
filter5[6][384] = 35'b11111011011100101100011010100000000;
filter5[6][385] = 35'b00000010101110010010011101001100000;
filter5[6][386] = 35'b00000100110101010101011101111000000;
filter5[6][387] = 35'b00000001101010011110001000010000000;
filter5[6][388] = 35'b00000001111110100111111110110100000;
filter5[6][389] = 35'b00000011010110001011010010101000000;
filter5[6][390] = 35'b00000010100111000001100101110000000;
filter5[6][391] = 35'b11111110110000001011011100100010000;
filter5[6][392] = 35'b11111110101100010001011101110100000;
filter5[6][393] = 35'b00000001101111001100011100001000000;
filter5[6][394] = 35'b00000001111010010011010000000000000;
filter5[6][395] = 35'b11111110110001001101110101100010000;
filter5[6][396] = 35'b11111110110010111001111001010000000;
filter5[6][397] = 35'b00000010101111100100111000011100000;
filter5[6][398] = 35'b00000101011111010111011001111000000;
filter5[6][399] = 35'b11111111111010100000100000111001100;
filter5[6][400] = 35'b11111100010001001111110110101000000;
filter5[6][401] = 35'b00000001100000010001110010100000000;
filter5[6][402] = 35'b11111111001110111000010110000101000;
filter5[6][403] = 35'b11111110101011111011011010110110000;
filter5[6][404] = 35'b11111111001110010001110001111000000;
filter5[6][405] = 35'b11111111011001111111000111001101000;
filter5[6][406] = 35'b11111111111110101101000001000000010;
filter5[6][407] = 35'b00000001110000001111110001010100000;
filter5[6][408] = 35'b00000000000000100011110010101000000;
filter5[6][409] = 35'b00000000010111100100110110000101100;
filter5[6][410] = 35'b11111010010111101010111000100000000;
filter5[6][411] = 35'b11111111010001110100100000110010000;
filter5[6][412] = 35'b00000000101001100001100001100001000;
filter5[6][413] = 35'b11111111101101001010010000000100000;
filter5[6][414] = 35'b00000101011100000111111000111000000;
filter5[6][415] = 35'b00000110101010001001101100011000000;
filter5[6][416] = 35'b00000010000011010010100010111100000;
filter5[6][417] = 35'b11111101111101110001001100100100000;
filter5[6][418] = 35'b00000010001111110110011110010100000;
filter5[6][419] = 35'b11111110001101001000100101101100000;
filter5[6][420] = 35'b00000000000011010001110100100101100;
filter5[6][421] = 35'b11111110001111000000100000101110000;
filter5[6][422] = 35'b11111110111000011000001111011100000;
filter5[6][423] = 35'b11111110111000110101001110100000000;
filter5[6][424] = 35'b11111101110011010110000011010100000;
filter5[6][425] = 35'b00000000010101010000010101000001000;
filter5[6][426] = 35'b00000000011010000110001001011111000;
filter5[6][427] = 35'b00000001001100101111010011100110000;
filter5[6][428] = 35'b11111110010101000000010101101100000;
filter5[6][429] = 35'b11110110110001100110111010110000000;
filter5[6][430] = 35'b11111101000110010000110101110100000;
filter5[6][431] = 35'b00000001000101011000010001111010000;
filter5[6][432] = 35'b11111111011111110011011000001100000;
filter5[6][433] = 35'b11111101100101011110001011101100000;
filter5[6][434] = 35'b11111111010000011000010000011110000;
filter5[6][435] = 35'b00000000111100000110000100010110000;
filter5[6][436] = 35'b11111101110101110101100000000100000;
filter5[6][437] = 35'b11111100011101000100110011010000000;
filter5[6][438] = 35'b11111110100010100001100001001010000;
filter5[6][439] = 35'b00000000000100000100001011111100111;
filter5[6][440] = 35'b11111111110111000001110110001001010;
filter5[6][441] = 35'b00000100110110101110000001111000000;
filter5[6][442] = 35'b11111101011011111001101100000000000;
filter5[6][443] = 35'b00000001101011111001111011100010000;
filter5[6][444] = 35'b00000011001000110111110101101100000;
filter5[6][445] = 35'b11111111001111110111000001010111000;
filter5[6][446] = 35'b11111101001010111010011010110000000;
filter5[6][447] = 35'b11111000101010111100000110111000000;
filter5[6][448] = 35'b11111111100110010100010110100011100;
filter5[6][449] = 35'b00000010101101001111110000101000000;
filter5[6][450] = 35'b00000100010010001010001010110000000;
filter5[6][451] = 35'b11111101001000001100110110010100000;
filter5[6][452] = 35'b00000011001100000001111001110000000;
filter5[6][453] = 35'b11111110010010010010110100001000000;
filter5[6][454] = 35'b11111111101111111111011111110011100;
filter5[6][455] = 35'b00000011011110100111000000100100000;
filter5[6][456] = 35'b00000001011110100100110101111000000;
filter5[6][457] = 35'b00000100001101100001111010011000000;
filter5[6][458] = 35'b11110111110010111010111100110000000;
filter5[6][459] = 35'b11111111110001011000000101111101000;
filter5[6][460] = 35'b11111111111101001101110101100001010;
filter5[6][461] = 35'b11110110001111110001101111010000000;
filter5[6][462] = 35'b11111111010010111000110010110000000;
filter5[6][463] = 35'b11111010100011010100001001100000000;
filter5[6][464] = 35'b11111110111010110001011100111100000;
filter5[6][465] = 35'b00000001100111100000010110011110000;
filter5[6][466] = 35'b11111110000111100010101100100010000;
filter5[6][467] = 35'b11111010111010000011010011010000000;
filter5[6][468] = 35'b11101111111001000010001110000000000;
filter5[6][469] = 35'b11110111100011000101100110110000000;
filter5[6][470] = 35'b11111000111000101011010111100000000;
filter5[6][471] = 35'b00000100100001001001100011011000000;
filter5[6][472] = 35'b00001001110111011001010111110000000;
filter5[6][473] = 35'b00000010000010101111001011010000000;
filter5[6][474] = 35'b00001010100101010010100001010000000;
filter5[6][475] = 35'b00000011101110110101110001100000000;
filter5[6][476] = 35'b11111010110110111001000010010000000;
filter5[6][477] = 35'b11111000100000010000101000101000000;
filter5[6][478] = 35'b11110110010100101010000001010000000;
filter5[6][479] = 35'b11111011010001100101101001000000000;
filter5[6][480] = 35'b00000001011010000111101011101000000;
filter5[6][481] = 35'b11111101110101011010111001001000000;
filter5[6][482] = 35'b00000001110000011110001001000000000;
filter5[6][483] = 35'b11111111100110101100010110001000000;
filter5[6][484] = 35'b11111000100100110011101010100000000;
filter5[6][485] = 35'b11111000100001101001001101001000000;
filter5[6][486] = 35'b11111111010000001011111010100111000;
filter5[6][487] = 35'b00000011110011100001000011100100000;
filter5[6][488] = 35'b11110101001110111110101010100000000;
filter5[6][489] = 35'b11111110001111111010001101110010000;
filter5[6][490] = 35'b00000000011100101011000101100110100;
filter5[6][491] = 35'b11111111100011111010011100000111000;
filter5[6][492] = 35'b11111001111000101011011101000000000;
filter5[6][493] = 35'b11111110101001001111010011000010000;
filter5[6][494] = 35'b00000000001001111111100010011011100;
filter5[6][495] = 35'b00000100001101110101010100110000000;
filter5[6][496] = 35'b11111110111111110100110000101000000;
filter5[6][497] = 35'b11111010101110010100001011001000000;
filter5[6][498] = 35'b11111110001011110110101111101110000;
filter5[6][499] = 35'b11111100110011001001111011100100000;
filter5[6][500] = 35'b00000001110010110000011011011100000;
filter5[6][501] = 35'b00000011111001000110110101011000000;
filter5[6][502] = 35'b11111111010101000010100011011001000;
filter5[6][503] = 35'b00000100010011010101101100100000000;
filter5[6][504] = 35'b00000001010110010110000010110110000;
filter5[6][505] = 35'b00000100110010111110000111001000000;
filter5[6][506] = 35'b11111001111000111000100100000000000;
filter5[6][507] = 35'b00000010100110000111000110111100000;
filter5[6][508] = 35'b00000000110101001001011101010001000;
filter5[6][509] = 35'b00000010000011010000000111001100000;
filter5[6][510] = 35'b11111011100001100111011000110000000;
filter5[6][511] = 35'b00000111100001101111101100110000000;
filter5[6][512] = 35'b00000100011000011100000001111000000;
filter5[6][513] = 35'b00000000010111001001001101111101000;
filter5[6][514] = 35'b00000001100101111110100000100110000;
filter5[6][515] = 35'b00000000001011010101011100111001110;
filter5[6][516] = 35'b00000010101000001100111101010000000;
filter5[6][517] = 35'b00000111001011000101001100100000000;
filter5[6][518] = 35'b00000000110000101011100011000001000;
filter5[6][519] = 35'b00000000100001100001011001000011000;
filter5[6][520] = 35'b11111110010100010110000011100110000;
filter5[6][521] = 35'b00000000011101010001110010111111100;
filter5[6][522] = 35'b00000011100010000000010110000100000;
filter5[6][523] = 35'b11111100111101101011001000011100000;
filter5[6][524] = 35'b00000001010100111010100000000100000;
filter5[6][525] = 35'b00000011000101111101000010000000000;
filter5[6][526] = 35'b00000010011001000101101111000000000;
filter5[6][527] = 35'b00000000000100000000100001001100111;
filter5[6][528] = 35'b11111101111001011010100010000100000;
filter5[6][529] = 35'b00000000001011000101000000011111100;
filter5[6][530] = 35'b11111100110111101000110111011100000;
filter5[6][531] = 35'b11111101011100000001011010011000000;
filter5[6][532] = 35'b00000001001001011010010100100100000;
filter5[6][533] = 35'b00000000011110100010110011101000000;
filter5[6][534] = 35'b11111110010001011011001000111100000;
filter5[6][535] = 35'b00000010110001011000111111001000000;
filter5[6][536] = 35'b11111110001001101001101111000110000;
filter5[6][537] = 35'b00000010010011110101111110001000000;
filter5[6][538] = 35'b11111101011100110001000001011000000;
filter5[6][539] = 35'b11111011011100010000001000001000000;
filter5[6][540] = 35'b00000001010111011101000011001010000;
filter5[6][541] = 35'b11111111111101010001001101011111011;
filter5[6][542] = 35'b00000010111111011100111010110100000;
filter5[6][543] = 35'b00000000101010011110001000100100000;
filter5[6][544] = 35'b11111111111010111001011111101010000;
filter5[6][545] = 35'b11111101011111101111111010110000000;
filter5[6][546] = 35'b00000000010011010010000110101111100;
filter5[6][547] = 35'b00000011100111110101110011101000000;
filter5[6][548] = 35'b11111110001101000001111110101010000;
filter5[6][549] = 35'b11111110010010000101111111101010000;
filter5[6][550] = 35'b11111110101011001001011101011100000;
filter5[6][551] = 35'b11111111100100101010111010011101000;
filter5[6][552] = 35'b11111001011110100110001100000000000;
filter5[6][553] = 35'b00000000110011111101001010110101000;
filter5[6][554] = 35'b11111110001111001111010100111110000;
filter5[6][555] = 35'b11111010010011100101100110110000000;
filter5[6][556] = 35'b11111101111000100011011111111100000;
filter5[6][557] = 35'b11111110011010011101011010111110000;
filter5[6][558] = 35'b11111010101110110111110110110000000;
filter5[6][559] = 35'b00000001110001110101110111100000000;
filter5[6][560] = 35'b11111100010110000000101011011100000;
filter5[6][561] = 35'b00000010100010011001100101100100000;
filter5[6][562] = 35'b00000010101010010110001010101100000;
filter5[6][563] = 35'b11111101001001001000011111110100000;
filter5[6][564] = 35'b00000001001100101000101010000110000;
filter5[6][565] = 35'b00000011000110010010011001010000000;
filter5[6][566] = 35'b00000100100101001110001011011000000;
filter5[6][567] = 35'b11111110110100110110001011001110000;
filter5[6][568] = 35'b11111001001011010000101111010000000;
filter5[6][569] = 35'b00000001111001001100010111011110000;
filter5[6][570] = 35'b00000000100011110000000010110101000;
filter5[6][571] = 35'b11111100100010110111011110000000000;
filter5[6][572] = 35'b00000010101101101111111010111000000;
filter5[6][573] = 35'b00000011000111010100001000101000000;
filter5[6][574] = 35'b00000010001001001110101001001100000;
filter5[6][575] = 35'b00000010110011010100011011001000000;
filter5[6][576] = 35'b00000000111011111110110111110100000;
filter5[6][577] = 35'b00000001010110011100110011010110000;
filter5[6][578] = 35'b00000011000110110011011011001000000;
filter5[6][579] = 35'b11111111110010000101001101110010000;
filter5[6][580] = 35'b00000000010000110010101101010101100;
filter5[6][581] = 35'b00000010011100010100100100001000000;
filter5[6][582] = 35'b00000011001011111011001001110000000;
filter5[6][583] = 35'b00000001000100011101111000001100000;
filter5[6][584] = 35'b11111000000111111110000001110000000;
filter5[6][585] = 35'b00000000011011001011100010001100000;
filter5[6][586] = 35'b11111101101000011001000110101000000;
filter5[6][587] = 35'b11111001110111010101110011110000000;
filter5[6][588] = 35'b00000000100001111111000010100111000;
filter5[6][589] = 35'b00000110101111011111010000011000000;
filter5[6][590] = 35'b00000110010101100110111100111000000;
filter5[6][591] = 35'b11111111001010011010000000001101000;
filter5[6][592] = 35'b11111101001110101011010001001100000;
filter5[6][593] = 35'b00000010000110111010010100001000000;
filter5[6][594] = 35'b11111011010101001011011110010000000;
filter5[6][595] = 35'b00000001011011100001101000110100000;
filter5[6][596] = 35'b11111101110101111000000011111100000;
filter5[6][597] = 35'b00000001101110100001111001100010000;
filter5[6][598] = 35'b00000001110001011110110110100110000;
filter5[6][599] = 35'b00000000011011000101101111011111000;
filter5[6][600] = 35'b11111110000010110001001000100010000;
filter5[6][601] = 35'b00000000001100110111000100010111000;
filter5[6][602] = 35'b11111110101110111001001000010010000;
filter5[6][603] = 35'b11111110010010001101100011101100000;
filter5[6][604] = 35'b00000000011001110110010001011001000;
filter5[6][605] = 35'b00000010000011010010010010001100000;
filter5[6][606] = 35'b00000010001101111100111110111000000;
filter5[6][607] = 35'b00000001100100011101111001101010000;
filter5[6][608] = 35'b00000001111000010110001000111110000;
filter5[6][609] = 35'b00000000111111000010001111000100000;
filter5[6][610] = 35'b11111110010111100110101000101100000;
filter5[6][611] = 35'b00000000000000110110001001001011101;
filter5[6][612] = 35'b11111011011100100000101010101000000;
filter5[6][613] = 35'b11111111101110000111110010101011000;
filter5[6][614] = 35'b11111101110001010000111010010100000;
filter5[6][615] = 35'b11111110110110110111011101001000000;
filter5[6][616] = 35'b00000000000010001100111101110100110;
filter5[6][617] = 35'b11111111011110111101001011111000000;
filter5[6][618] = 35'b11111011000111001001101111011000000;
filter5[6][619] = 35'b11111101101101000111000101110000000;
filter5[6][620] = 35'b00000001001001100011011110110010000;
filter5[6][621] = 35'b00000010101001110111001101111100000;
filter5[6][622] = 35'b11111011101110001010110111100000000;
filter5[6][623] = 35'b11111110110010110101110111010110000;
filter5[6][624] = 35'b11111100101110001101111010010000000;
filter5[6][625] = 35'b00000010100101001011011000001100000;
filter5[6][626] = 35'b11110110110100001000011000010000000;
filter5[6][627] = 35'b11111011001101001100000000000000000;
filter5[6][628] = 35'b00000000010110111000010111100101000;
filter5[6][629] = 35'b00000101011110110101010001001000000;
filter5[6][630] = 35'b00000010010001101111011101110100000;
filter5[6][631] = 35'b11111111011110110011111000101111000;
filter5[6][632] = 35'b00000001010011010101001101001000000;
filter5[6][633] = 35'b00000011101100110101010110110100000;
filter5[6][634] = 35'b11110110011101110111011100010000000;
filter5[6][635] = 35'b11111010011100001011011100100000000;
filter5[6][636] = 35'b00000000000011100111110010101101111;
filter5[6][637] = 35'b00000010001001011110011001101000000;
filter5[6][638] = 35'b00000011000001111101011110001000000;
filter5[6][639] = 35'b00000101001001001110100011010000000;
filter5[6][640] = 35'b11111110101111101000000100101110000;
filter5[6][641] = 35'b00000011010111010011100001110100000;
filter5[6][642] = 35'b00001010010101000011011010110000000;
filter5[6][643] = 35'b11111110000000010101001110011110000;
filter5[6][644] = 35'b11111111011010110111000111111010000;
filter5[6][645] = 35'b11111111001011101111011000010011000;
filter5[6][646] = 35'b11111100100001000010000111111100000;
filter5[6][647] = 35'b11111000110111111010011010000000000;
filter5[6][648] = 35'b11111110010000101000110111100000000;
filter5[6][649] = 35'b00000011110111110010100000001100000;
filter5[6][650] = 35'b00000000110100101000100010000111000;
filter5[6][651] = 35'b11111101111010001110111010111100000;
filter5[6][652] = 35'b00000011011001100111011111000000000;
filter5[6][653] = 35'b11111111110001100101000100001010110;
filter5[6][654] = 35'b11111110010110100010100001001010000;
filter5[6][655] = 35'b11111010010101110001111110110000000;
filter5[6][656] = 35'b00000010011101000101110001000100000;
filter5[6][657] = 35'b00000011010100100000000000100000000;
filter5[6][658] = 35'b00000000000100001110110011110110100;
filter5[6][659] = 35'b00000000001101010100110000000010100;
filter5[6][660] = 35'b11111011100000010100110111101000000;
filter5[6][661] = 35'b00000010000101110011101011111000000;
filter5[6][662] = 35'b00000110011011100001011010001000000;
filter5[6][663] = 35'b00000101010010111011100000000000000;
filter5[6][664] = 35'b00000010001111110110001100111000000;
filter5[6][665] = 35'b11111110100101111001101000110010000;
filter5[6][666] = 35'b11111010011001010011101100001000000;
filter5[6][667] = 35'b11111111001100111010010101000110000;
filter5[6][668] = 35'b11111111100111011001110010010010100;
filter5[6][669] = 35'b00000010100110001110000011000000000;
filter5[6][670] = 35'b00000100101001010101111010000000000;
filter5[6][671] = 35'b00000010101101000111010111101000000;
filter5[6][672] = 35'b11111101110000101010110001110100000;
filter5[6][673] = 35'b11111011101001010111110001101000000;
filter5[6][674] = 35'b11111011100100110000010101110000000;
filter5[6][675] = 35'b11111100011011111010000010010000000;
filter5[6][676] = 35'b11111010011111101101111010110000000;
filter5[6][677] = 35'b00000000101110001100111101101010000;
filter5[6][678] = 35'b11111110010010001001100110010110000;
filter5[6][679] = 35'b00000011010010011110110000100000000;
filter5[6][680] = 35'b11110100101111110011011100010000000;
filter5[6][681] = 35'b11111110110001010100001010000010000;
filter5[6][682] = 35'b00000010010101011110011001110000000;
filter5[6][683] = 35'b11111100101110100110010110110100000;
filter5[6][684] = 35'b11111000100000111111000101011000000;
filter5[6][685] = 35'b11111111111111000111100011011110011;
filter5[6][686] = 35'b11111100000101011101001100101100000;
filter5[6][687] = 35'b00001000000111001001011001100000000;
filter5[6][688] = 35'b11111001011010101101111101110000000;
filter5[6][689] = 35'b11111111111100110010101100100101000;
filter5[6][690] = 35'b00000001101110101001010100101010000;
filter5[6][691] = 35'b00000000111010000101110110010100000;
filter5[6][692] = 35'b11111101101001011000111010001000000;
filter5[6][693] = 35'b00000001011011010011001101000100000;
filter5[6][694] = 35'b11111110101100010101000011111000000;
filter5[6][695] = 35'b00000010010010100111001011010000000;
filter5[6][696] = 35'b00000000011011110001101011011011100;
filter5[6][697] = 35'b00000000001000100010111010001001010;
filter5[6][698] = 35'b11111101001110001110100010111000000;
filter5[6][699] = 35'b00000000011110010101101010001111000;
filter5[6][700] = 35'b00000010001101100101100111011100000;
filter5[6][701] = 35'b00000000000110001110001001110001010;
filter5[6][702] = 35'b11111101101110110010000111110100000;
filter5[6][703] = 35'b11111011100100010000111111000000000;
filter5[6][704] = 35'b11111100001011000101111111101100000;
filter5[6][705] = 35'b11111111000000011100000001111010000;
filter5[6][706] = 35'b11111101101110101001100110100100000;
filter5[6][707] = 35'b11111100001011010110011101010100000;
filter5[6][708] = 35'b11111111011001101001110101101101000;
filter5[6][709] = 35'b11111111000101101110011001111010000;
filter5[6][710] = 35'b00000001111101010101100001001110000;
filter5[6][711] = 35'b11111101000010001010000110010000000;
filter5[6][712] = 35'b00000000001000100011111010011100000;
filter5[6][713] = 35'b11111110000111011110010111001100000;
filter5[6][714] = 35'b11111100011100101001100110001100000;
filter5[6][715] = 35'b11111111110110000100000111001010110;
filter5[6][716] = 35'b11111100011110010111111001100000000;
filter5[6][717] = 35'b00000001111101001000011001010010000;
filter5[6][718] = 35'b11111101101110010111011011101100000;
filter5[6][719] = 35'b00000000010110011001111000111011100;
filter5[6][720] = 35'b11111110011010101101101011101010000;
filter5[6][721] = 35'b11111100010010010101111011010100000;
filter5[6][722] = 35'b00000000000101111010101111000111100;
filter5[6][723] = 35'b00000000010100011001001011001100100;
filter5[6][724] = 35'b00000001100110101101010111010110000;
filter5[6][725] = 35'b00000000001011100111001000101101100;
filter5[6][726] = 35'b00000001001000000001111000010100000;
filter5[6][727] = 35'b00000000000010011110010111101011000;
filter5[6][728] = 35'b11111111110111000110001001111111000;
filter5[6][729] = 35'b11111011101001110001001001100000000;
filter5[6][730] = 35'b11111110110000111100110111110010000;
filter5[6][731] = 35'b11111111100011000010010011001100000;
filter5[6][732] = 35'b00000010001101010100000011001000000;
filter5[6][733] = 35'b11111111110111101010001110001010110;
filter5[6][734] = 35'b11111101111011010100001101010000000;
filter5[6][735] = 35'b11111110100010010100011000111110000;
filter5[6][736] = 35'b11111010011101010101111111100000000;
filter5[6][737] = 35'b11111010011011101111110101100000000;
filter5[6][738] = 35'b00000001101110111110011111100010000;
filter5[6][739] = 35'b00000000101001100111101111101000000;
filter5[6][740] = 35'b11111110001010000101101000011100000;
filter5[6][741] = 35'b11111111010000100110100111010010000;
filter5[6][742] = 35'b11111100111010010101110111011000000;
filter5[6][743] = 35'b00000000001100000110011111010111110;
filter5[6][744] = 35'b11111101000001000011001100001100000;
filter5[6][745] = 35'b00000001010011010001011011101000000;
filter5[6][746] = 35'b11111011101000011101001010000000000;
filter5[6][747] = 35'b11111111011000001011110000110100000;
filter5[6][748] = 35'b11111110101010000001111100000100000;
filter5[6][749] = 35'b00000010101010010010101100011100000;
filter5[6][750] = 35'b00000000100011110010111100011101000;
filter5[6][751] = 35'b00000001001100001000110100100100000;
filter5[6][752] = 35'b11111111010110010110001100011101000;
filter5[6][753] = 35'b11111111100101011011000001110001100;
filter5[6][754] = 35'b11111100010100111101101010110000000;
filter5[6][755] = 35'b11111011010001001111100111101000000;
filter5[6][756] = 35'b00000001111110010101111100010010000;
filter5[6][757] = 35'b00000010000110111011110101011100000;
filter5[6][758] = 35'b00000010110011100110000011000100000;
filter5[6][759] = 35'b00000100010100100001000110111000000;
filter5[6][760] = 35'b11111100110101001110011010110100000;
filter5[6][761] = 35'b00000000000011110110111010000100000;
filter5[6][762] = 35'b11111010111101001101000010100000000;
filter5[6][763] = 35'b11111101101111110100000111010000000;
filter5[6][764] = 35'b00000110010110100010111000111000000;
filter5[6][765] = 35'b00000101010010101011101010101000000;
filter5[6][766] = 35'b00000001011001000111101001110110000;
filter5[6][767] = 35'b00000011100001010111111111110100000;
filter5[6][768] = 35'b00000100110010110110001011010000000;
filter5[6][769] = 35'b00000100110000101010010110101000000;
filter5[6][770] = 35'b11111110100111110010101001000010000;
filter5[6][771] = 35'b00000011000011110011111010111100000;
filter5[6][772] = 35'b00000101011111001110111101011000000;
filter5[6][773] = 35'b00000100000000101011001001010000000;
filter5[6][774] = 35'b11111010111001100110100100010000000;
filter5[6][775] = 35'b11111111011110001001001011011100000;
filter5[6][776] = 35'b00000000000001101011000010000010111;
filter5[6][777] = 35'b00000011001000010100001111001100000;
filter5[6][778] = 35'b00000110110100010101111010011000000;
filter5[6][779] = 35'b11111101011111100100111000100000000;
filter5[6][780] = 35'b11111111101101110000000010001111100;
filter5[6][781] = 35'b00000000110001100001101100100011000;
filter5[6][782] = 35'b11111101011111001101101001011000000;
filter5[6][783] = 35'b00000010111001101001110011111000000;
filter5[6][784] = 35'b00000000111101001100010010010010000;
filter5[6][785] = 35'b00000011001100000000100100011100000;
filter5[6][786] = 35'b00000011100000011101110010010000000;
filter5[6][787] = 35'b00000000101101111011000101101000000;
filter5[6][788] = 35'b11111110110100000100101010000100000;
filter5[6][789] = 35'b11111100000011111101001010100100000;
filter5[6][790] = 35'b00000000101010011100011110000101000;
filter5[6][791] = 35'b11111100111111011010110001010000000;
filter5[6][792] = 35'b00000000100101101000010101010110000;
filter5[6][793] = 35'b00000011000011100100101001100100000;
filter5[6][794] = 35'b00000100010001010110011010010000000;
filter5[6][795] = 35'b11111011001101111010111100101000000;
filter5[6][796] = 35'b11111110010010111100011111111000000;
filter5[6][797] = 35'b11111000100010111100110100011000000;
filter5[6][798] = 35'b11111011101011111110101000111000000;
filter5[6][799] = 35'b11111101010010010101001101100100000;
filter5[6][800] = 35'b11111101101010111110100010100000000;
filter5[6][801] = 35'b00000001101111101000100010000000000;
filter5[6][802] = 35'b00000000110000110101001110011101000;
filter5[6][803] = 35'b11111110001111110111011110100110000;
filter5[6][804] = 35'b11111101101110000011110100010000000;
filter5[6][805] = 35'b11110101101101101010100100000000000;
filter5[6][806] = 35'b11111001001100001111001110011000000;
filter5[6][807] = 35'b11111111110010100110101000110010010;
filter5[6][808] = 35'b11111111010011001100000111010010000;
filter5[6][809] = 35'b11111100011111010010111011010000000;
filter5[6][810] = 35'b11111011110101110100010001001000000;
filter5[6][811] = 35'b11111011001000100100011001001000000;
filter5[6][812] = 35'b11111011111010100010111011001000000;
filter5[6][813] = 35'b11111110010001101100100010100100000;
filter5[6][814] = 35'b00000001101010100101000101010000000;
filter5[6][815] = 35'b00000100011011001001100001010000000;
filter5[6][816] = 35'b11111111101101000101000100000011000;
filter5[6][817] = 35'b00000000011011101000111011110000100;
filter5[6][818] = 35'b00000000010111000001000000010011000;
filter5[6][819] = 35'b11111101101100000100000000101000000;
filter5[6][820] = 35'b11111001001110101111000010101000000;
filter5[6][821] = 35'b00000011000101110101011111010100000;
filter5[6][822] = 35'b00000010000011101100110000100000000;
filter5[6][823] = 35'b00000110111111111101011110011000000;
filter5[6][824] = 35'b00000000011010011001111111100010100;
filter5[6][825] = 35'b00000000111100000011100000101010000;
filter5[6][826] = 35'b00000011001001000001010111110000000;
filter5[6][827] = 35'b11111110000110101000011011010010000;
filter5[6][828] = 35'b11111100011011111001100111100000000;
filter5[6][829] = 35'b00000011110111000010110000101000000;
filter5[6][830] = 35'b11111110110110000111101111000110000;
filter5[6][831] = 35'b00000111101111011000000000011000000;
filter5[6][832] = 35'b11111110001010000001000110110100000;
filter5[6][833] = 35'b11111101101000000100101000100100000;
filter5[6][834] = 35'b11111011111000101110000000001000000;
filter5[6][835] = 35'b11111101100111111110100111101100000;
filter5[6][836] = 35'b11111101110000010100101110010000000;
filter5[6][837] = 35'b11111110001111011101111001111110000;
filter5[6][838] = 35'b11111101011000111000011011001000000;
filter5[6][839] = 35'b11111110101010011100101010001010000;
filter5[6][840] = 35'b11111101101000100000010111111000000;
filter5[6][841] = 35'b11111111011100001001110001010000000;
filter5[6][842] = 35'b11111011110011010001011110010000000;
filter5[6][843] = 35'b11111111000000000011100101010110000;
filter5[6][844] = 35'b00000001011010000101001001011100000;
filter5[6][845] = 35'b11111110100010110000100000010100000;
filter5[6][846] = 35'b00000000101000001100111111101101000;
filter5[6][847] = 35'b11111110010110110010100001110000000;
filter5[6][848] = 35'b11111111001110101111011001010101000;
filter5[6][849] = 35'b11111101101110000111101101100100000;
filter5[6][850] = 35'b11111101101010000001001011010100000;
filter5[6][851] = 35'b11111011101010100111010100011000000;
filter5[6][852] = 35'b00000011001001101101001101000000000;
filter5[6][853] = 35'b00000010100101100111000100101100000;
filter5[6][854] = 35'b00000001011110111101101111110100000;
filter5[6][855] = 35'b11111110101000011110110011000000000;
filter5[6][856] = 35'b00000000001110001101111110011101000;
filter5[6][857] = 35'b11111010101010000100111011000000000;
filter5[6][858] = 35'b11111011111100101110010000011000000;
filter5[6][859] = 35'b00000001110010011111010110010010000;
filter5[6][860] = 35'b00000001110110101100000010010100000;
filter5[6][861] = 35'b00000001000101100101010101011110000;
filter5[6][862] = 35'b11111011011101000110000111111000000;
filter5[6][863] = 35'b11111010000111111000101111110000000;
filter5[6][864] = 35'b11111111100011111001011011000000100;
filter5[6][865] = 35'b11111100110010110011110111100000000;
filter5[6][866] = 35'b00000010010010001011101010101100000;
filter5[6][867] = 35'b11111111110011101010101001001111110;
filter5[6][868] = 35'b00000010111110110001000111010100000;
filter5[6][869] = 35'b00000000000010111111101010000000010;
filter5[6][870] = 35'b11111101000000101100100100111000000;
filter5[6][871] = 35'b00000010001010111100010011010100000;
filter5[6][872] = 35'b11111010110111111100010111001000000;
filter5[6][873] = 35'b11111110011100110010110110110010000;
filter5[6][874] = 35'b11111101111111000010100111100100000;
filter5[6][875] = 35'b00000010101101100001000001101100000;
filter5[6][876] = 35'b11111110110111111010110111111000000;
filter5[6][877] = 35'b00000000110110100110011101100011000;
filter5[6][878] = 35'b00000010101101011011010001000100000;
filter5[6][879] = 35'b11111111001001110001111101001100000;
filter5[6][880] = 35'b11111101110110111110010001110000000;
filter5[6][881] = 35'b00000000001001101010101111001001100;
filter5[6][882] = 35'b11111010010000001101100110101000000;
filter5[6][883] = 35'b11111101101100010000111111011000000;
filter5[6][884] = 35'b00000010010111110111110100011000000;
filter5[6][885] = 35'b00000100000011111101111100011000000;
filter5[6][886] = 35'b00000011001010011101001110111000000;
filter5[6][887] = 35'b00000000010001111000100010011011100;
filter5[6][888] = 35'b11111100010001110001110011011000000;
filter5[6][889] = 35'b11111111101111101001000010001101000;
filter5[6][890] = 35'b11111010001101000001010111001000000;
filter5[6][891] = 35'b11111011110111101111001110010000000;
filter5[6][892] = 35'b00000010101011111111000011100100000;
filter5[6][893] = 35'b11111101000010110011110111110100000;
filter5[6][894] = 35'b00001001011101001001000111100000000;
filter5[6][895] = 35'b11111110110101100000111000010000000;
filter5[6][896] = 35'b11110101001100110101100100010000000;
filter5[6][897] = 35'b11111111101000101001111100001111000;
filter5[6][898] = 35'b11111000111111100101100001000000000;
filter5[6][899] = 35'b11110111110011110111010000110000000;
filter5[6][900] = 35'b11111111000101001000110001101001000;
filter5[6][901] = 35'b00000101110010100011100110101000000;
filter5[6][902] = 35'b00000001011111001111100100111100000;
filter5[6][903] = 35'b11111001110001111011111011110000000;
filter5[6][904] = 35'b11110111001110011000100010000000000;
filter5[6][905] = 35'b11110011010001101000011100100000000;
filter5[6][906] = 35'b11110000001010011000001111110000000;
filter5[6][907] = 35'b00000001111010101010101011111110000;
filter5[6][908] = 35'b00000000101101111011000010011110000;
filter5[6][909] = 35'b00000000111100111010011000101100000;
filter5[6][910] = 35'b11111110101101111010001001111000000;
filter5[6][911] = 35'b00001000000000011101111000100000000;
filter5[6][912] = 35'b00000010101110101000110000010100000;
filter5[6][913] = 35'b11101110100001101000101010100000000;
filter5[6][914] = 35'b11111100010100100000101011010100000;
filter5[6][915] = 35'b00000001011100010000111010100100000;
filter5[6][916] = 35'b00000000010101100011100000101001100;
filter5[6][917] = 35'b11111111010001101010101101100100000;
filter5[6][918] = 35'b00000000000011000101010110111001011;
filter5[6][919] = 35'b11111111001000011011101100111111000;
filter5[6][920] = 35'b11111010000001110000100101001000000;
filter5[6][921] = 35'b11110111101101101000101010110000000;
filter5[6][922] = 35'b11111101110100101100011100010100000;
filter5[6][923] = 35'b00000010011111001111001100110100000;
filter5[6][924] = 35'b00000001001010010001111100100000000;
filter5[6][925] = 35'b00000000010000101000101001001001000;
filter5[6][926] = 35'b11111101110110011001101000110000000;
filter5[6][927] = 35'b00000001000100000100100111110000000;
filter5[6][928] = 35'b11111001001011101000010010000000000;
filter5[6][929] = 35'b11111111101001110101100010101011100;
filter5[6][930] = 35'b00000011010000001001101110011100000;
filter5[6][931] = 35'b11111111010101011101111001110101000;
filter5[6][932] = 35'b00000000101011001101001010110110000;
filter5[6][933] = 35'b11111111011101011010011101100111000;
filter5[6][934] = 35'b11111100100100111110000110110100000;
filter5[6][935] = 35'b00000100111001001011111000100000000;
filter5[6][936] = 35'b00000001101110011011111110011110000;
filter5[6][937] = 35'b00000000000011100110110101101011100;
filter5[6][938] = 35'b11111111101101101111001111001011000;
filter5[6][939] = 35'b11111101001111100100010101001100000;
filter5[6][940] = 35'b00000010001111111000010100100100000;
filter5[6][941] = 35'b00000011001011110100110101101100000;
filter5[6][942] = 35'b00000010001000011100111010111000000;
filter5[6][943] = 35'b00000011101001101001000011100000000;
filter5[6][944] = 35'b00000000100100010100011110001011000;
filter5[6][945] = 35'b00000010010111101111110100110100000;
filter5[6][946] = 35'b11111101011001110101010111010000000;
filter5[6][947] = 35'b11111010010001011001001000010000000;
filter5[6][948] = 35'b00000011111011101001011001010100000;
filter5[6][949] = 35'b00000000101101101011001000110110000;
filter5[6][950] = 35'b11111010001001001100101100100000000;
filter5[6][951] = 35'b00000011011010001101011000001100000;
filter5[6][952] = 35'b11111110011010100101000001111100000;
filter5[6][953] = 35'b11110010000101110100011000100000000;
filter5[6][954] = 35'b00000001101010011000100110100110000;
filter5[6][955] = 35'b00000000101010101101100110100011000;
filter5[6][956] = 35'b00000000001011011100001111010000100;
filter5[6][957] = 35'b00000100000110110011000001000000000;
filter5[6][958] = 35'b00001000100100100001010110010000000;
filter5[6][959] = 35'b00000001100000011110110010011010000;
filter5[6][960] = 35'b00000000010101001110111011000110000;
filter5[6][961] = 35'b11111110101000011000010000110010000;
filter5[6][962] = 35'b11111101101001111010101011110100000;
filter5[6][963] = 35'b11110101110001100111111001000000000;
filter5[6][964] = 35'b11111111010001000111000011111110000;
filter5[6][965] = 35'b00000011101100110011101101110100000;
filter5[6][966] = 35'b00000110100001110111101101110000000;
filter5[6][967] = 35'b00000011011111101010000110010000000;
filter5[6][968] = 35'b11111110110101111111110001101010000;
filter5[6][969] = 35'b11111100010001100110000001011100000;
filter5[6][970] = 35'b11111011001001000010101010101000000;
filter5[6][971] = 35'b00000010000000100101001101101100000;
filter5[6][972] = 35'b11111101001101011011100011000000000;
filter5[6][973] = 35'b00000000011111100000011110010001000;
filter5[6][974] = 35'b00000010001110100111100011001000000;
filter5[6][975] = 35'b00000000111101001101000000010001000;
filter5[6][976] = 35'b11110111010100101001111001000000000;
filter5[6][977] = 35'b11110101010111100100010101100000000;
filter5[6][978] = 35'b00000001110101110110100010010100000;
filter5[6][979] = 35'b00000010100111011110011100010100000;
filter5[6][980] = 35'b11111110000110101110001011111110000;
filter5[6][981] = 35'b00000000001110111110101111011111100;
filter5[6][982] = 35'b00000001100000110010111011001000000;
filter5[6][983] = 35'b00000001100100000001111101101110000;
filter5[6][984] = 35'b11110011111101011100100100000000000;
filter5[6][985] = 35'b11111101011011101010100010010100000;
filter5[6][986] = 35'b00000010010010110001010001101000000;
filter5[6][987] = 35'b00000111001000011010010001001000000;
filter5[6][988] = 35'b11111110011011111010110100101110000;
filter5[6][989] = 35'b11111010011010000001110111010000000;
filter5[6][990] = 35'b11111111111101111001110101100000111;
filter5[6][991] = 35'b00000001001101011011101101100110000;
filter5[6][992] = 35'b11111011000011101000100100010000000;
filter5[6][993] = 35'b11110111101110001000010110100000000;
filter5[6][994] = 35'b11110111101001001000111110100000000;
filter5[6][995] = 35'b11111111000110101111011110111101000;
filter5[6][996] = 35'b00000000101011001101011100101010000;
filter5[6][997] = 35'b00000001110100101001100111110100000;
filter5[6][998] = 35'b00000010100110000100100100111100000;
filter5[6][999] = 35'b11111001011110110100101101101000000;
filter5[6][1000] = 35'b11111100000000011000100100100100000;
filter5[6][1001] = 35'b11111100100000100101010110100100000;
filter5[6][1002] = 35'b11110100100111010100101101100000000;
filter5[6][1003] = 35'b11111000110000011111011111000000000;
filter5[6][1004] = 35'b00000010010100110110100010010000000;
filter5[6][1005] = 35'b00000010110010101001001111000000000;
filter5[6][1006] = 35'b11111110001111011011001101110100000;
filter5[6][1007] = 35'b00000010110111111111111110001000000;
filter5[6][1008] = 35'b11111101001010010100001101000100000;
filter5[6][1009] = 35'b11111101010101101011110010110100000;
filter5[6][1010] = 35'b11110000100100000011101110010000000;
filter5[6][1011] = 35'b11111000110111001001100010000000000;
filter5[6][1012] = 35'b00000000110001000011000000111010000;
filter5[6][1013] = 35'b00000111001000001001011011010000000;
filter5[6][1014] = 35'b00001001111011100101111100110000000;
filter5[6][1015] = 35'b11111101101101100001100001101100000;
filter5[6][1016] = 35'b11111011001000011111000111001000000;
filter5[6][1017] = 35'b11111001100001001000001110010000000;
filter5[6][1018] = 35'b11111010011010100001100101000000000;
filter5[6][1019] = 35'b00000101110110001011001010110000000;
filter5[6][1020] = 35'b00000111100000101001100110010000000;
filter5[6][1021] = 35'b00000010001000101011100011001000000;
filter5[6][1022] = 35'b00000111010111101000101011101000000;
filter5[6][1023] = 35'b11111101000000001101010100000000000;
filter5[7][0] = 35'b11111111101111010101111000110011000;
filter5[7][1] = 35'b11111101011101000100011000001000000;
filter5[7][2] = 35'b11111101111000000101100100000100000;
filter5[7][3] = 35'b00000000100011011000011001111110000;
filter5[7][4] = 35'b00000010100011111110000111001100000;
filter5[7][5] = 35'b00000011000101101101110110011100000;
filter5[7][6] = 35'b00000000000010101011100001100001000;
filter5[7][7] = 35'b00000010111101000100111110101100000;
filter5[7][8] = 35'b00000000111000000010011010110011000;
filter5[7][9] = 35'b00000101101111001100111111010000000;
filter5[7][10] = 35'b00001010000010100010000111100000000;
filter5[7][11] = 35'b11111110111100011011011111101010000;
filter5[7][12] = 35'b11111110000001001011110011110000000;
filter5[7][13] = 35'b00000010011011101010001111011100000;
filter5[7][14] = 35'b00000110000011100110001101011000000;
filter5[7][15] = 35'b11111101110011100000000000101100000;
filter5[7][16] = 35'b11111111000000111101101111101001000;
filter5[7][17] = 35'b00000010110000100000011001110100000;
filter5[7][18] = 35'b00000100110000000101100100011000000;
filter5[7][19] = 35'b00000000110110101001010100010111000;
filter5[7][20] = 35'b00000001110101001010011001000000000;
filter5[7][21] = 35'b00000001100100000100110111100000000;
filter5[7][22] = 35'b00000011101101100100101001111100000;
filter5[7][23] = 35'b00000010001011110011000010000100000;
filter5[7][24] = 35'b11111011101001110001110100111000000;
filter5[7][25] = 35'b11111100010010011110001010011000000;
filter5[7][26] = 35'b00000001000010110110110111001000000;
filter5[7][27] = 35'b00000000010011001000100000001101100;
filter5[7][28] = 35'b00000010101001110110100011100100000;
filter5[7][29] = 35'b11111111010100101110010100101111000;
filter5[7][30] = 35'b00000010100111010000100001111100000;
filter5[7][31] = 35'b11111110000011100111010111001010000;
filter5[7][32] = 35'b00000001011111011011101110100110000;
filter5[7][33] = 35'b11111110100011011000101011110100000;
filter5[7][34] = 35'b11111011001011010111100000001000000;
filter5[7][35] = 35'b11111111011111011010010001011011000;
filter5[7][36] = 35'b00000000001010011110100101110110010;
filter5[7][37] = 35'b11110100111011101000110001110000000;
filter5[7][38] = 35'b11110011110110101110111011010000000;
filter5[7][39] = 35'b00000101010011010011110111011000000;
filter5[7][40] = 35'b00000000100101010011010011001010000;
filter5[7][41] = 35'b00000000101110001100010110010101000;
filter5[7][42] = 35'b00000001010110111101001111011110000;
filter5[7][43] = 35'b00000001000001111010111011101010000;
filter5[7][44] = 35'b11111010001110011100110101001000000;
filter5[7][45] = 35'b11111000101011011110100101011000000;
filter5[7][46] = 35'b11110010100100001000001001000000000;
filter5[7][47] = 35'b00000011111011110000101100001100000;
filter5[7][48] = 35'b00000001001101111101100111000110000;
filter5[7][49] = 35'b00000000000100001011111000010001011;
filter5[7][50] = 35'b11111101101101111010010100001000000;
filter5[7][51] = 35'b00000111101100001001110011001000000;
filter5[7][52] = 35'b11110100010111110010111000100000000;
filter5[7][53] = 35'b11101100111010010111011111100000000;
filter5[7][54] = 35'b00000010000000001110001111010100000;
filter5[7][55] = 35'b00000011100100111011101010100000000;
filter5[7][56] = 35'b11111110111100011100011110101000000;
filter5[7][57] = 35'b00000101101010111010110100010000000;
filter5[7][58] = 35'b11111110001111110010110110010100000;
filter5[7][59] = 35'b00000101100001001101011000100000000;
filter5[7][60] = 35'b11111010010000111011111100100000000;
filter5[7][61] = 35'b00000001011000101001001011001110000;
filter5[7][62] = 35'b00000101111011101111111110101000000;
filter5[7][63] = 35'b00001010010001111001000110100000000;
filter5[7][64] = 35'b00000000111100111001100111110000000;
filter5[7][65] = 35'b00000010011111110100000010010000000;
filter5[7][66] = 35'b11111100111101101111011001011100000;
filter5[7][67] = 35'b00000010101111011101100100101000000;
filter5[7][68] = 35'b00000011000001101101010101010000000;
filter5[7][69] = 35'b11111111000110110000100111100110000;
filter5[7][70] = 35'b11111100011101011110001011001000000;
filter5[7][71] = 35'b11111101001110000000111110001100000;
filter5[7][72] = 35'b11111100000010001010001100000100000;
filter5[7][73] = 35'b11111111110110110000011101000001000;
filter5[7][74] = 35'b00000110101110000101110011110000000;
filter5[7][75] = 35'b11111010111110011100100001100000000;
filter5[7][76] = 35'b00000011001101000011000111111100000;
filter5[7][77] = 35'b00000011001111001000110001111000000;
filter5[7][78] = 35'b00000000000010110010111000000111101;
filter5[7][79] = 35'b00000011010110010101100011110100000;
filter5[7][80] = 35'b11111110110101101011001110100110000;
filter5[7][81] = 35'b00000001001100010111111111000100000;
filter5[7][82] = 35'b00000010010101101010011010111000000;
filter5[7][83] = 35'b11111110111011110001110011000110000;
filter5[7][84] = 35'b11111111100101101101001000010010100;
filter5[7][85] = 35'b00000001010110111101010001110100000;
filter5[7][86] = 35'b11111100000111110001000011011000000;
filter5[7][87] = 35'b00000010010001100010001101000000000;
filter5[7][88] = 35'b11111100001001111001111010011100000;
filter5[7][89] = 35'b11110111111101101001000001110000000;
filter5[7][90] = 35'b11111111011010011101010111011111000;
filter5[7][91] = 35'b00000001001100110101111111110110000;
filter5[7][92] = 35'b00000010110010000101011111001100000;
filter5[7][93] = 35'b00000000110100011110011001110011000;
filter5[7][94] = 35'b11111101010110110001100110001000000;
filter5[7][95] = 35'b11111011000000010111100010011000000;
filter5[7][96] = 35'b11111111110110010000101101001110010;
filter5[7][97] = 35'b11111101111111111001100100011000000;
filter5[7][98] = 35'b11111011101111101011011110001000000;
filter5[7][99] = 35'b11111111011101110110011101100101000;
filter5[7][100] = 35'b11111111010000100111110101101101000;
filter5[7][101] = 35'b11111111001101101011010101101011000;
filter5[7][102] = 35'b00000011010010010101000111111000000;
filter5[7][103] = 35'b11111101100100100001010011010100000;
filter5[7][104] = 35'b11111111011010111111111110000001000;
filter5[7][105] = 35'b00000001101001111110100111101100000;
filter5[7][106] = 35'b00000001011100011111101100011110000;
filter5[7][107] = 35'b11111110000001100111111111000100000;
filter5[7][108] = 35'b11111011111110111100010011110000000;
filter5[7][109] = 35'b00000000011110110111011100010000100;
filter5[7][110] = 35'b00000011010100010001110100110000000;
filter5[7][111] = 35'b11111110010101111001111010100010000;
filter5[7][112] = 35'b00000001101101011110011110010000000;
filter5[7][113] = 35'b11111110100000011101100001010100000;
filter5[7][114] = 35'b11111111101010110101100001000010000;
filter5[7][115] = 35'b00000001001110010010110110111000000;
filter5[7][116] = 35'b00000000111101110001010111110101000;
filter5[7][117] = 35'b11111100100011101110101111010000000;
filter5[7][118] = 35'b00000110010101000111000111100000000;
filter5[7][119] = 35'b00000001101010101010111110100100000;
filter5[7][120] = 35'b00000100000000101100000010010000000;
filter5[7][121] = 35'b11111101101000011001011100010000000;
filter5[7][122] = 35'b11111101011101101011101010100100000;
filter5[7][123] = 35'b00000011010011101111011011100000000;
filter5[7][124] = 35'b00000010110100011000100110000100000;
filter5[7][125] = 35'b00000000001110100001011010001010110;
filter5[7][126] = 35'b11111011000010111110110001011000000;
filter5[7][127] = 35'b00000001111000110101100110001100000;
filter5[7][128] = 35'b11110111011010110111100100110000000;
filter5[7][129] = 35'b00000001001010001010110100001110000;
filter5[7][130] = 35'b11110110101010010111110101010000000;
filter5[7][131] = 35'b11111101011101100010110011000000000;
filter5[7][132] = 35'b11101111000010000011001110100000000;
filter5[7][133] = 35'b11110101010011111000110000010000000;
filter5[7][134] = 35'b11111000100101101001100000111000000;
filter5[7][135] = 35'b11111011111111100001011000011000000;
filter5[7][136] = 35'b00000100010001001101110010101000000;
filter5[7][137] = 35'b00000000001101100101010100010000010;
filter5[7][138] = 35'b11110011111001111010000101100000000;
filter5[7][139] = 35'b11101000010010000010010100100000000;
filter5[7][140] = 35'b00000000001010100011011010110011110;
filter5[7][141] = 35'b11110100000110100011001100100000000;
filter5[7][142] = 35'b11101010000001111011100101100000000;
filter5[7][143] = 35'b11111001101001001010000001101000000;
filter5[7][144] = 35'b11111010101000001101110111111000000;
filter5[7][145] = 35'b11110010001111110011110010110000000;
filter5[7][146] = 35'b11110100000111100010011111000000000;
filter5[7][147] = 35'b11111110001010101001011001010110000;
filter5[7][148] = 35'b11111101011110010001001111111000000;
filter5[7][149] = 35'b00000010001011111001000110000100000;
filter5[7][150] = 35'b11101100110011111001001011000000000;
filter5[7][151] = 35'b11110110000100011100000110100000000;
filter5[7][152] = 35'b11110110100011110011101100100000000;
filter5[7][153] = 35'b11110111011100011000101101100000000;
filter5[7][154] = 35'b11111100111111101101101100110100000;
filter5[7][155] = 35'b00000000100101011010001100101000000;
filter5[7][156] = 35'b00000010100010010100101111100000000;
filter5[7][157] = 35'b00000000100101110001110011010010000;
filter5[7][158] = 35'b11110111001001100000011011110000000;
filter5[7][159] = 35'b11111010111100010110000111111000000;
filter5[7][160] = 35'b11110010100010010101001011110000000;
filter5[7][161] = 35'b11111100101000111101001111111000000;
filter5[7][162] = 35'b00000010100000011111111001100100000;
filter5[7][163] = 35'b00000001011101101010100100111010000;
filter5[7][164] = 35'b00000001000011101001101110011000000;
filter5[7][165] = 35'b11111110110001110101111000000100000;
filter5[7][166] = 35'b00000011010111001110001101010100000;
filter5[7][167] = 35'b11110001001101110111010000110000000;
filter5[7][168] = 35'b11111111111000111110001100011100111;
filter5[7][169] = 35'b11111110110001101000101011101000000;
filter5[7][170] = 35'b00000110101101001100110111110000000;
filter5[7][171] = 35'b11111111000101001001110001110110000;
filter5[7][172] = 35'b11111101010111101100110011100100000;
filter5[7][173] = 35'b11111101011100101010111100010000000;
filter5[7][174] = 35'b00000001110111011010011111011100000;
filter5[7][175] = 35'b11111011000100001110001110111000000;
filter5[7][176] = 35'b00000111001101111001100111100000000;
filter5[7][177] = 35'b00001001000001001110001001100000000;
filter5[7][178] = 35'b00001110010101000100101001010000000;
filter5[7][179] = 35'b00000100010000001011001011001000000;
filter5[7][180] = 35'b11111011110011111101110011100000000;
filter5[7][181] = 35'b00000010101100111110110110001000000;
filter5[7][182] = 35'b11111111010011010100111101000000000;
filter5[7][183] = 35'b11101010101000001110000101100000000;
filter5[7][184] = 35'b00000101001110100000110001010000000;
filter5[7][185] = 35'b00000001100001111111000001101110000;
filter5[7][186] = 35'b11111011111111001100100100011000000;
filter5[7][187] = 35'b11111001000111001001001000111000000;
filter5[7][188] = 35'b11111011011011100110111101100000000;
filter5[7][189] = 35'b00001011011110000101100010010000000;
filter5[7][190] = 35'b11111101001111110001100000111000000;
filter5[7][191] = 35'b11110111010010001010100001010000000;
filter5[7][192] = 35'b11111100100011001011101001110100000;
filter5[7][193] = 35'b11101100001010100110111100000000000;
filter5[7][194] = 35'b00000011111001010011101110101000000;
filter5[7][195] = 35'b00000101010000001000011111000000000;
filter5[7][196] = 35'b00000110101011010111011101100000000;
filter5[7][197] = 35'b00000101010101101011000110111000000;
filter5[7][198] = 35'b00000001011111110110011001011010000;
filter5[7][199] = 35'b11111101010010011010011011011100000;
filter5[7][200] = 35'b00000100010101101000001100011000000;
filter5[7][201] = 35'b11111010100110011011001110111000000;
filter5[7][202] = 35'b11111000101111100101011011001000000;
filter5[7][203] = 35'b00000011101110011100100001011000000;
filter5[7][204] = 35'b11111001010111001001111011010000000;
filter5[7][205] = 35'b11110111101101101101010010000000000;
filter5[7][206] = 35'b00000110101110101010010011111000000;
filter5[7][207] = 35'b00000001000001001111100010001010000;
filter5[7][208] = 35'b11111101110101101100111000000000000;
filter5[7][209] = 35'b11111010110001100011110101100000000;
filter5[7][210] = 35'b11111011110101010000001110101000000;
filter5[7][211] = 35'b00000011101010100001011010011000000;
filter5[7][212] = 35'b00000011110000101000000110000000000;
filter5[7][213] = 35'b00000101001000010010110101000000000;
filter5[7][214] = 35'b11111011110100011010001110000000000;
filter5[7][215] = 35'b11101100111010111110110001100000000;
filter5[7][216] = 35'b11110011111010010111111001100000000;
filter5[7][217] = 35'b00000101100010010101111001000000000;
filter5[7][218] = 35'b11101010101000101110111011000000000;
filter5[7][219] = 35'b11111110111110101001111011100000000;
filter5[7][220] = 35'b00000000010000001110100100111001000;
filter5[7][221] = 35'b11111011110011100001101110011000000;
filter5[7][222] = 35'b11110110111101011111100001110000000;
filter5[7][223] = 35'b00000110011111111100010010110000000;
filter5[7][224] = 35'b11111000000011110100010110000000000;
filter5[7][225] = 35'b11111111100101111011110001001010100;
filter5[7][226] = 35'b00000100100011110001111010110000000;
filter5[7][227] = 35'b11111010000010000101110110100000000;
filter5[7][228] = 35'b00000001111101010011111110011000000;
filter5[7][229] = 35'b11111101110100111101000011101000000;
filter5[7][230] = 35'b11111100111110101110011100110100000;
filter5[7][231] = 35'b11110101111101000001010101100000000;
filter5[7][232] = 35'b11111011110111110001010111101000000;
filter5[7][233] = 35'b11111110101001001010111010000110000;
filter5[7][234] = 35'b00000010011110110100110111110100000;
filter5[7][235] = 35'b11111100010001010010100110100100000;
filter5[7][236] = 35'b00000001100101100101110011001010000;
filter5[7][237] = 35'b00000000111001110001001110111001000;
filter5[7][238] = 35'b00000100001101011100100101100000000;
filter5[7][239] = 35'b11111000010100110010000010100000000;
filter5[7][240] = 35'b00000000111111010111110110100001000;
filter5[7][241] = 35'b00000100010000110000001111110000000;
filter5[7][242] = 35'b00000000100010000100010100000011000;
filter5[7][243] = 35'b11111111100111101001100000110000100;
filter5[7][244] = 35'b11111111011011000100111100001110000;
filter5[7][245] = 35'b00000001110110010001101100001000000;
filter5[7][246] = 35'b11111111101010001111001010100011100;
filter5[7][247] = 35'b00000010000101011101011110100000000;
filter5[7][248] = 35'b11111011010010100101000001111000000;
filter5[7][249] = 35'b00000101111101100011000000110000000;
filter5[7][250] = 35'b11111100111010000110110111110000000;
filter5[7][251] = 35'b11111110111010100000110010010010000;
filter5[7][252] = 35'b00000001110111111101110100010110000;
filter5[7][253] = 35'b11111110111011000101110010001000000;
filter5[7][254] = 35'b11110110110110110101110010110000000;
filter5[7][255] = 35'b11111010001011000001110001111000000;
filter5[7][256] = 35'b11111101010000100000100001111000000;
filter5[7][257] = 35'b11111100101100111110011101001100000;
filter5[7][258] = 35'b00000011011111111110111100110100000;
filter5[7][259] = 35'b00000000101101110000010011011101000;
filter5[7][260] = 35'b00000000110110000100010001010100000;
filter5[7][261] = 35'b11111111101111000110101100110111100;
filter5[7][262] = 35'b00000001100111100011000111010000000;
filter5[7][263] = 35'b11111111000101101110001011100010000;
filter5[7][264] = 35'b11111111111110001111111001011010101;
filter5[7][265] = 35'b11111100000001100111010110001000000;
filter5[7][266] = 35'b11111100101011100011100000001000000;
filter5[7][267] = 35'b11111001001011111111010100010000000;
filter5[7][268] = 35'b11111000000010011100100011100000000;
filter5[7][269] = 35'b11111000001000111011011111111000000;
filter5[7][270] = 35'b00000001010100100010001111111000000;
filter5[7][271] = 35'b00000111100000000011011111111000000;
filter5[7][272] = 35'b11111000010110110100100111001000000;
filter5[7][273] = 35'b11101101011011100100001011100000000;
filter5[7][274] = 35'b11100111100100101111010001100000000;
filter5[7][275] = 35'b00000111110101101011010000101000000;
filter5[7][276] = 35'b00000001101011111100001001110100000;
filter5[7][277] = 35'b11110111010010100011110101110000000;
filter5[7][278] = 35'b11110001100010100011100111100000000;
filter5[7][279] = 35'b11111101011110111111101001110100000;
filter5[7][280] = 35'b11110011010000101011110001110000000;
filter5[7][281] = 35'b11110110010100010101001010000000000;
filter5[7][282] = 35'b00000001111001001100101101011100000;
filter5[7][283] = 35'b11111001011011111110011110001000000;
filter5[7][284] = 35'b11111001100011010001001010100000000;
filter5[7][285] = 35'b11111111111101101000111111001000001;
filter5[7][286] = 35'b11110100110101111000111100110000000;
filter5[7][287] = 35'b11110101111100001011101010110000000;
filter5[7][288] = 35'b11110100010100000011100011000000000;
filter5[7][289] = 35'b11110010111001001011001100100000000;
filter5[7][290] = 35'b00000010010000010001101000000000000;
filter5[7][291] = 35'b00000001110010100111011000001010000;
filter5[7][292] = 35'b11111111110111000110001101001110010;
filter5[7][293] = 35'b00000100110000110010100000111000000;
filter5[7][294] = 35'b11111101101000110111011111000100000;
filter5[7][295] = 35'b11110100110000101011011000010000000;
filter5[7][296] = 35'b11111101100010100011110010001000000;
filter5[7][297] = 35'b11110001010100111001100001000000000;
filter5[7][298] = 35'b00000001000010000010011110001110000;
filter5[7][299] = 35'b11111110111111111110011100100100000;
filter5[7][300] = 35'b00000010011100110001000001101000000;
filter5[7][301] = 35'b00000001001100111101001101000010000;
filter5[7][302] = 35'b11111111110100100011000111100101100;
filter5[7][303] = 35'b11111001110101111010001110111000000;
filter5[7][304] = 35'b00001010010011001100110111100000000;
filter5[7][305] = 35'b00000000000110101111001000101101110;
filter5[7][306] = 35'b11111101011001001110111101001000000;
filter5[7][307] = 35'b00000011110100001101011101010100000;
filter5[7][308] = 35'b11111110110011010100010000111100000;
filter5[7][309] = 35'b11111110011010001010010001101100000;
filter5[7][310] = 35'b11111011110010110101010110000000000;
filter5[7][311] = 35'b11110111000010011001101011110000000;
filter5[7][312] = 35'b11111100011001101110101010101000000;
filter5[7][313] = 35'b11110010011100001000100111000000000;
filter5[7][314] = 35'b00000000000110111001110100000101101;
filter5[7][315] = 35'b00000000101110110011000010001101000;
filter5[7][316] = 35'b11111100101001110110010000101100000;
filter5[7][317] = 35'b00000001000110110111001111001010000;
filter5[7][318] = 35'b11110110010100000110100101110000000;
filter5[7][319] = 35'b11110100011111110111011011010000000;
filter5[7][320] = 35'b00000000011001110100000111101110100;
filter5[7][321] = 35'b11111111100111110000000110011001000;
filter5[7][322] = 35'b00000100000100001000101101100000000;
filter5[7][323] = 35'b11111111101110111001001000110111000;
filter5[7][324] = 35'b00000110110110001010010101000000000;
filter5[7][325] = 35'b11111011010111100111101000001000000;
filter5[7][326] = 35'b11111101111110001110001000100000000;
filter5[7][327] = 35'b00000100101001111101011101010000000;
filter5[7][328] = 35'b11111111001011110001011010110101000;
filter5[7][329] = 35'b00000011001001001101000100100100000;
filter5[7][330] = 35'b00000000011100101000100001001101100;
filter5[7][331] = 35'b00000000101000010101100110100000000;
filter5[7][332] = 35'b11111101111111100100110010110100000;
filter5[7][333] = 35'b11111110011100101011010100010010000;
filter5[7][334] = 35'b00000000101101011000110010011001000;
filter5[7][335] = 35'b11111101100111100000010011110100000;
filter5[7][336] = 35'b00000000100101101101111001010001000;
filter5[7][337] = 35'b00000000100100000010011000000111000;
filter5[7][338] = 35'b11111110001011010001000110111100000;
filter5[7][339] = 35'b11111111011101110111110110010010000;
filter5[7][340] = 35'b00000001001100111100100110011110000;
filter5[7][341] = 35'b00000100101111010110110110000000000;
filter5[7][342] = 35'b00000011111100101111000101000100000;
filter5[7][343] = 35'b11111111000010010110101010110111000;
filter5[7][344] = 35'b11111001000110100101111010001000000;
filter5[7][345] = 35'b11111111000001011111001000010001000;
filter5[7][346] = 35'b11111100110000000000001011101000000;
filter5[7][347] = 35'b11111111000001101101000010100001000;
filter5[7][348] = 35'b00000010111110110000010111011100000;
filter5[7][349] = 35'b11111100000100110001001000000100000;
filter5[7][350] = 35'b11110111110010111000001101000000000;
filter5[7][351] = 35'b11111110101101101110100101101110000;
filter5[7][352] = 35'b11111111111000101110111000010011010;
filter5[7][353] = 35'b11111110111111011101011100001000000;
filter5[7][354] = 35'b00000000001001010110100001011001010;
filter5[7][355] = 35'b11111111000111011010100010000101000;
filter5[7][356] = 35'b00000010001101010000000011010100000;
filter5[7][357] = 35'b11111010001111101101100101100000000;
filter5[7][358] = 35'b00000000110110010000010110000000000;
filter5[7][359] = 35'b11111111000111111101111001001101000;
filter5[7][360] = 35'b11111110010100100111010001010110000;
filter5[7][361] = 35'b00000010111010000010001110110000000;
filter5[7][362] = 35'b00001000000000100010111010100000000;
filter5[7][363] = 35'b11111110100111101100001011101100000;
filter5[7][364] = 35'b11111100111100010011111100011000000;
filter5[7][365] = 35'b11111111000010101101010110111010000;
filter5[7][366] = 35'b00000011111011111011001011111100000;
filter5[7][367] = 35'b11111111100000001011111010101111000;
filter5[7][368] = 35'b11111110010010010111011001010000000;
filter5[7][369] = 35'b00000100000100010101000101000000000;
filter5[7][370] = 35'b11111011001001110011001110111000000;
filter5[7][371] = 35'b11111101101111111011011110110000000;
filter5[7][372] = 35'b00000001010101101100010111010110000;
filter5[7][373] = 35'b11111110110010011111001100010010000;
filter5[7][374] = 35'b11111111101010101111001001000011100;
filter5[7][375] = 35'b11111111000111000110010001101101000;
filter5[7][376] = 35'b00000001011011001001110010010100000;
filter5[7][377] = 35'b00000100000101110110000101011000000;
filter5[7][378] = 35'b11110111010010000001010101000000000;
filter5[7][379] = 35'b00000001100010000000101101110110000;
filter5[7][380] = 35'b00000011111100101110111010000100000;
filter5[7][381] = 35'b11111011110000011010101011011000000;
filter5[7][382] = 35'b11111010000001100110110100000000000;
filter5[7][383] = 35'b00000001000001100111001110010110000;
filter5[7][384] = 35'b11111110100111011000011111011110000;
filter5[7][385] = 35'b00000000100100011010111011110101000;
filter5[7][386] = 35'b11111111010101101110100111110000000;
filter5[7][387] = 35'b11111111111000001000001001101110001;
filter5[7][388] = 35'b00000000010010000111010000000011100;
filter5[7][389] = 35'b00000000101010101110110101001100000;
filter5[7][390] = 35'b00000000001001101010010000011100110;
filter5[7][391] = 35'b00000001110111000010111011111000000;
filter5[7][392] = 35'b11111101110001101101101111010100000;
filter5[7][393] = 35'b00000001101000110001001101000100000;
filter5[7][394] = 35'b00000010101101110011011100000000000;
filter5[7][395] = 35'b00000000010110010110010001110110000;
filter5[7][396] = 35'b11111110000110001111111110100000000;
filter5[7][397] = 35'b11111101011100110101100110111100000;
filter5[7][398] = 35'b00000100010010011110000001110000000;
filter5[7][399] = 35'b00000001111101011111011100011000000;
filter5[7][400] = 35'b11111110000101110100000101011110000;
filter5[7][401] = 35'b11111101101011000010111011010100000;
filter5[7][402] = 35'b00000001111011101110111010010000000;
filter5[7][403] = 35'b00000000001110111110001110001010100;
filter5[7][404] = 35'b11111101100101111000010100101000000;
filter5[7][405] = 35'b00000001101100100101000100011000000;
filter5[7][406] = 35'b00000011101011110010101111001100000;
filter5[7][407] = 35'b00000001000001100101100001011000000;
filter5[7][408] = 35'b11111011011110111010001110000000000;
filter5[7][409] = 35'b11111101101011001110011000100000000;
filter5[7][410] = 35'b00000001011010110001110011100110000;
filter5[7][411] = 35'b11111110111101101001000000110100000;
filter5[7][412] = 35'b00000000011110101111011011000000000;
filter5[7][413] = 35'b11111110111010001011110011001100000;
filter5[7][414] = 35'b11111111111110010110101010101000110;
filter5[7][415] = 35'b11111111101111010110000001001101000;
filter5[7][416] = 35'b11111100011111100101110000000000000;
filter5[7][417] = 35'b11111110001111100101100110110010000;
filter5[7][418] = 35'b11111101110111110000110101110000000;
filter5[7][419] = 35'b11111101101010101000001000101100000;
filter5[7][420] = 35'b11111111001001000001000011110011000;
filter5[7][421] = 35'b00000001011110110100001100000010000;
filter5[7][422] = 35'b00000000101011100101001110001011000;
filter5[7][423] = 35'b00000001110011111110011011001000000;
filter5[7][424] = 35'b11111110110001100011110001111100000;
filter5[7][425] = 35'b00000001001001011000000111111100000;
filter5[7][426] = 35'b00000001111110010101000110000000000;
filter5[7][427] = 35'b11111100011100011101000011001000000;
filter5[7][428] = 35'b11111100011100000000101011111100000;
filter5[7][429] = 35'b00000000100011101101111110110110000;
filter5[7][430] = 35'b11111100011100000111001001110100000;
filter5[7][431] = 35'b00000001110100010100101110010010000;
filter5[7][432] = 35'b00000000100001000010101001010101000;
filter5[7][433] = 35'b00000011100001101010100011101000000;
filter5[7][434] = 35'b11111100111110001111110001000100000;
filter5[7][435] = 35'b11110110110010110011110010100000000;
filter5[7][436] = 35'b11111100010100100100001111111100000;
filter5[7][437] = 35'b11111110000101110000000000001100000;
filter5[7][438] = 35'b00000100101101001111101100000000000;
filter5[7][439] = 35'b00000001001111111101001101001000000;
filter5[7][440] = 35'b11111111110010000111111110100000110;
filter5[7][441] = 35'b11111111101101011110000101011111000;
filter5[7][442] = 35'b11111111011110111000111011101110000;
filter5[7][443] = 35'b11111100111111011001100110000000000;
filter5[7][444] = 35'b11111111001001011011011111001101000;
filter5[7][445] = 35'b00000001001001110000001101111100000;
filter5[7][446] = 35'b11111110100100101001011000010100000;
filter5[7][447] = 35'b00000001011111000001100010101000000;
filter5[7][448] = 35'b11111111111100100111011100000101101;
filter5[7][449] = 35'b11111010001111011101101101111000000;
filter5[7][450] = 35'b11111100110000000011000110100000000;
filter5[7][451] = 35'b00000010000011001101000001101100000;
filter5[7][452] = 35'b00000001001000000101101111101000000;
filter5[7][453] = 35'b11111110000110001100100010010000000;
filter5[7][454] = 35'b00000010000001000000101001111000000;
filter5[7][455] = 35'b00000100000001111010011001000000000;
filter5[7][456] = 35'b11111101111011110111100011111100000;
filter5[7][457] = 35'b00000000101001100011011110010011000;
filter5[7][458] = 35'b11111111001101010000010101001001000;
filter5[7][459] = 35'b00000010000001000001001110001000000;
filter5[7][460] = 35'b11111111000011111011110111011000000;
filter5[7][461] = 35'b00000100111010001001110101100000000;
filter5[7][462] = 35'b00000101110001001000111100100000000;
filter5[7][463] = 35'b11111110001011100010001111110110000;
filter5[7][464] = 35'b11111101010110110100010000101000000;
filter5[7][465] = 35'b00000000011110111101110100101101100;
filter5[7][466] = 35'b00000001000011001010100111111000000;
filter5[7][467] = 35'b11111110101100000110101111101100000;
filter5[7][468] = 35'b00000000010010010011110001000101000;
filter5[7][469] = 35'b00000000011101110000100010000011100;
filter5[7][470] = 35'b11111010111111001111110011010000000;
filter5[7][471] = 35'b00000000010010111001110101011101000;
filter5[7][472] = 35'b11111100111000011001110011101100000;
filter5[7][473] = 35'b00000000110110001111100011010101000;
filter5[7][474] = 35'b00000010001010100011101000000000000;
filter5[7][475] = 35'b11111110001101011010010111001010000;
filter5[7][476] = 35'b00000010110010001100001010101000000;
filter5[7][477] = 35'b11111111101110101001111111010100000;
filter5[7][478] = 35'b11111101011000110110111000101000000;
filter5[7][479] = 35'b00000001100010000100111010011100000;
filter5[7][480] = 35'b11111100111101010011100010100100000;
filter5[7][481] = 35'b11111010101101000111101101111000000;
filter5[7][482] = 35'b00001001010001100110011111110000000;
filter5[7][483] = 35'b00000000101001001001100010000110000;
filter5[7][484] = 35'b00000000100110010010100101111011000;
filter5[7][485] = 35'b00000001000001011011010101101100000;
filter5[7][486] = 35'b11111000001111100010011101110000000;
filter5[7][487] = 35'b11110011110100100101110100110000000;
filter5[7][488] = 35'b11111111100011000100000011001101100;
filter5[7][489] = 35'b00000101001111011111010010011000000;
filter5[7][490] = 35'b00000110001001000010001100011000000;
filter5[7][491] = 35'b11111110011100010001000010011000000;
filter5[7][492] = 35'b11111101001001111111010001101100000;
filter5[7][493] = 35'b00000011111000101000100000011100000;
filter5[7][494] = 35'b11111111011110101000011111110101000;
filter5[7][495] = 35'b11111101000011101101011101000100000;
filter5[7][496] = 35'b11111101011010111010000110011100000;
filter5[7][497] = 35'b00000011000010100010100010001100000;
filter5[7][498] = 35'b00001000100000110100001101010000000;
filter5[7][499] = 35'b00000010100000101000111010101100000;
filter5[7][500] = 35'b11111010010010111001000011011000000;
filter5[7][501] = 35'b00000000101100101001110001010111000;
filter5[7][502] = 35'b11111110110000001000000111010010000;
filter5[7][503] = 35'b00000001110100110010011000100100000;
filter5[7][504] = 35'b00000011001110000010110000001000000;
filter5[7][505] = 35'b11111100111101111011000100000000000;
filter5[7][506] = 35'b00000010010010110101111111101000000;
filter5[7][507] = 35'b11111100100011011011100011001000000;
filter5[7][508] = 35'b11111111010101100011010100100110000;
filter5[7][509] = 35'b00000000111000100111111011001100000;
filter5[7][510] = 35'b11111110000010010101000011000010000;
filter5[7][511] = 35'b00000001010101011001011110100100000;
filter5[7][512] = 35'b11111111101011001011100010110000000;
filter5[7][513] = 35'b11111101011000100100001000001000000;
filter5[7][514] = 35'b11111111011001100011011110111010000;
filter5[7][515] = 35'b00000001011101111100101100101100000;
filter5[7][516] = 35'b00000100011010010111101001011000000;
filter5[7][517] = 35'b11111101000111100101000110110100000;
filter5[7][518] = 35'b00000000101000111110001111011100000;
filter5[7][519] = 35'b11111010000000101001100000010000000;
filter5[7][520] = 35'b11111111010000001110011011011001000;
filter5[7][521] = 35'b00000010100101111000100100111000000;
filter5[7][522] = 35'b00000011110010100011011011000000000;
filter5[7][523] = 35'b11111110100010010000110011110100000;
filter5[7][524] = 35'b11111110011110110111011110010000000;
filter5[7][525] = 35'b00000011101101000101111100101000000;
filter5[7][526] = 35'b00000011010001011010010111110000000;
filter5[7][527] = 35'b00000100000111100000001111111000000;
filter5[7][528] = 35'b11111101100110101110000010110100000;
filter5[7][529] = 35'b00000100011000000101100101001000000;
filter5[7][530] = 35'b11111110111100000001111100100000000;
filter5[7][531] = 35'b11111111000110110111100101101110000;
filter5[7][532] = 35'b11111110111011001010110011100000000;
filter5[7][533] = 35'b11111100110101110110011110001000000;
filter5[7][534] = 35'b00000001011010010101101110110000000;
filter5[7][535] = 35'b11111111101001000001001011111101000;
filter5[7][536] = 35'b11111100110011110001000100000100000;
filter5[7][537] = 35'b00000000110001011000100101010000000;
filter5[7][538] = 35'b11111111010101101011101000110010000;
filter5[7][539] = 35'b11111110000010101100011001110100000;
filter5[7][540] = 35'b11111111010011001101011001000101000;
filter5[7][541] = 35'b11111110000000010110101100011100000;
filter5[7][542] = 35'b11111110010011100000100011100100000;
filter5[7][543] = 35'b11111110010110001001001000101000000;
filter5[7][544] = 35'b11111100100011110111010001010000000;
filter5[7][545] = 35'b00000001010100111010000000011100000;
filter5[7][546] = 35'b11111111110111010010110011111101000;
filter5[7][547] = 35'b11111101010100001100100010100100000;
filter5[7][548] = 35'b00000011000001010110001111000000000;
filter5[7][549] = 35'b11111011101101000110001111111000000;
filter5[7][550] = 35'b00000011111011000011101110001100000;
filter5[7][551] = 35'b11111111001100001010001100111001000;
filter5[7][552] = 35'b11111110011101111110000100110100000;
filter5[7][553] = 35'b11111101111101001010100001111100000;
filter5[7][554] = 35'b00000000110101111101011000110100000;
filter5[7][555] = 35'b11110100111111010010101110000000000;
filter5[7][556] = 35'b00000000000101111101100111101101111;
filter5[7][557] = 35'b00000010000110001111000101110100000;
filter5[7][558] = 35'b00000000000000101000011100100101000;
filter5[7][559] = 35'b00000011101011001110001111000000000;
filter5[7][560] = 35'b11111110010001101000101000000000000;
filter5[7][561] = 35'b11111101100110101001100010101000000;
filter5[7][562] = 35'b00000001001000000110011100010000000;
filter5[7][563] = 35'b11110111101100000011001011010000000;
filter5[7][564] = 35'b00000110100101101000011001001000000;
filter5[7][565] = 35'b00000000010111011101111011101111100;
filter5[7][566] = 35'b00000010000111011110111101111000000;
filter5[7][567] = 35'b00000001010001011011000101100110000;
filter5[7][568] = 35'b00000000011001001110001101111011000;
filter5[7][569] = 35'b00000100110010110110000010011000000;
filter5[7][570] = 35'b11111000110110011111110010011000000;
filter5[7][571] = 35'b11111010100011100001001111101000000;
filter5[7][572] = 35'b00001001101101110010111110000000000;
filter5[7][573] = 35'b11111110101011010100010010100100000;
filter5[7][574] = 35'b00000100010011110010110111010000000;
filter5[7][575] = 35'b11111110101011110111100100011010000;
filter5[7][576] = 35'b11111111110010111100010100111010010;
filter5[7][577] = 35'b11111101111001101100001011100000000;
filter5[7][578] = 35'b00000001110100100101011000110100000;
filter5[7][579] = 35'b00000000000100001100001011000010110;
filter5[7][580] = 35'b00000011111001110111000110010000000;
filter5[7][581] = 35'b11111110110011111010101011111010000;
filter5[7][582] = 35'b00000000111110010111011011100111000;
filter5[7][583] = 35'b11111111110111111101010000011101000;
filter5[7][584] = 35'b11111111110100100110001011011111010;
filter5[7][585] = 35'b00000010001010000000011000001000000;
filter5[7][586] = 35'b00000000110100010110001111010000000;
filter5[7][587] = 35'b11111110010111011011101101001100000;
filter5[7][588] = 35'b11111101100101111110101111110100000;
filter5[7][589] = 35'b11111101111111010111011000010000000;
filter5[7][590] = 35'b11111111100100001010100010110010000;
filter5[7][591] = 35'b00000010010100001110001001100000000;
filter5[7][592] = 35'b00000000001101111010000011011111100;
filter5[7][593] = 35'b00000011101000101110001010000000000;
filter5[7][594] = 35'b11111101000010010110111100010100000;
filter5[7][595] = 35'b11111111011100101101100000010011000;
filter5[7][596] = 35'b11111111100001110000000001110000000;
filter5[7][597] = 35'b11111111001101011100111000011100000;
filter5[7][598] = 35'b00000001110101111011101001100010000;
filter5[7][599] = 35'b00000001011111000011010011010000000;
filter5[7][600] = 35'b11111100000001011000001011110100000;
filter5[7][601] = 35'b11111111110001010100010010001000100;
filter5[7][602] = 35'b11111111110001110111010001000111110;
filter5[7][603] = 35'b11111100001000101111111111101100000;
filter5[7][604] = 35'b00000010000101111010100010110000000;
filter5[7][605] = 35'b11111101100100111101111000000000000;
filter5[7][606] = 35'b11111011010100111000101111000000000;
filter5[7][607] = 35'b00000001010100001000101010010100000;
filter5[7][608] = 35'b11111101011010001010110000100100000;
filter5[7][609] = 35'b11111110101111111101011110100110000;
filter5[7][610] = 35'b00000000011011100101001000001100100;
filter5[7][611] = 35'b00000000101110100100000010001110000;
filter5[7][612] = 35'b00000000010010000110000110001100000;
filter5[7][613] = 35'b11111101101110011010111000111100000;
filter5[7][614] = 35'b00000010001101000011000000000100000;
filter5[7][615] = 35'b11111110101000100110010010000100000;
filter5[7][616] = 35'b00000010100110110101101001110000000;
filter5[7][617] = 35'b11111100011100010000010111000100000;
filter5[7][618] = 35'b00000010101011101010001111100100000;
filter5[7][619] = 35'b00000011010101000110110111100100000;
filter5[7][620] = 35'b11111001010011011011100110110000000;
filter5[7][621] = 35'b11111111111000000100011100010000000;
filter5[7][622] = 35'b00000010001110110011110000010100000;
filter5[7][623] = 35'b11111111000101000111110000010001000;
filter5[7][624] = 35'b11111110101010010110111111110110000;
filter5[7][625] = 35'b00000100000110001001101110100000000;
filter5[7][626] = 35'b00000100100000011001111010110000000;
filter5[7][627] = 35'b00000010100000001000011110000100000;
filter5[7][628] = 35'b11111011010111110100001000001000000;
filter5[7][629] = 35'b00000010010010000001011001100000000;
filter5[7][630] = 35'b00000010010111101011010010100000000;
filter5[7][631] = 35'b11111100100000111101011110110100000;
filter5[7][632] = 35'b11111011111101000000110100100000000;
filter5[7][633] = 35'b11110111111110000111011100010000000;
filter5[7][634] = 35'b11111110111010100110010111110000000;
filter5[7][635] = 35'b00000000101001000110111011001110000;
filter5[7][636] = 35'b11111111001111110111011010000111000;
filter5[7][637] = 35'b11111110111101010001011001011000000;
filter5[7][638] = 35'b11111011101000100111000001101000000;
filter5[7][639] = 35'b00000011101101001111000101000000000;
filter5[7][640] = 35'b00000010011010110010111000110100000;
filter5[7][641] = 35'b11111101000110000001110010101000000;
filter5[7][642] = 35'b11111001101100010100000000101000000;
filter5[7][643] = 35'b00000001101100010101101111110110000;
filter5[7][644] = 35'b00000011000010001011111010001100000;
filter5[7][645] = 35'b11111100100000111010101011100100000;
filter5[7][646] = 35'b11111101100101100100010110001000000;
filter5[7][647] = 35'b00000000001000011011011010100011010;
filter5[7][648] = 35'b00000001011010110001110000000000000;
filter5[7][649] = 35'b11111110011111101101101111110110000;
filter5[7][650] = 35'b00000000100101000001010011101000000;
filter5[7][651] = 35'b11111111100111011011000000001001000;
filter5[7][652] = 35'b11111101001000011001111100000100000;
filter5[7][653] = 35'b11111110100111001100111100010000000;
filter5[7][654] = 35'b00000000101010110111110101011110000;
filter5[7][655] = 35'b11111001101000110010000001000000000;
filter5[7][656] = 35'b11111111110001110010101100110000010;
filter5[7][657] = 35'b11111101000011011010011100000100000;
filter5[7][658] = 35'b00000100001111010111000111100000000;
filter5[7][659] = 35'b00000111111101001001110101110000000;
filter5[7][660] = 35'b11111110111000110101011000011100000;
filter5[7][661] = 35'b11111100111101000001010111100000000;
filter5[7][662] = 35'b11111111011010001001101101010110000;
filter5[7][663] = 35'b11111000100101101010011110111000000;
filter5[7][664] = 35'b11111100110000011101000000011100000;
filter5[7][665] = 35'b11111110100110010001011100101100000;
filter5[7][666] = 35'b00000011101101001000010001010000000;
filter5[7][667] = 35'b00000110000011010001000001010000000;
filter5[7][668] = 35'b00000001111000101000110111011110000;
filter5[7][669] = 35'b00000000010101100111100111110010100;
filter5[7][670] = 35'b00000010001011100011011001001000000;
filter5[7][671] = 35'b11111111100001110101111000001000000;
filter5[7][672] = 35'b11111010111011110010000100101000000;
filter5[7][673] = 35'b11111100111100101011011011110100000;
filter5[7][674] = 35'b11111101011110100001010010011000000;
filter5[7][675] = 35'b11110111110010011000100001110000000;
filter5[7][676] = 35'b11111111101010000100111000010001000;
filter5[7][677] = 35'b11111011010111000101111000001000000;
filter5[7][678] = 35'b11111110010101000000000011001100000;
filter5[7][679] = 35'b00000010101101100101010001111000000;
filter5[7][680] = 35'b11111101000111000111111001001000000;
filter5[7][681] = 35'b11111110100100001000011110100010000;
filter5[7][682] = 35'b11110001001111110111010101110000000;
filter5[7][683] = 35'b11110111101100011100011100010000000;
filter5[7][684] = 35'b11111111001001000100000101101000000;
filter5[7][685] = 35'b00000010001111010000101111001000000;
filter5[7][686] = 35'b11111110111101111101000001001000000;
filter5[7][687] = 35'b00000010011010001011110000000100000;
filter5[7][688] = 35'b11111100100010010000111101001100000;
filter5[7][689] = 35'b00000000001000111000101100011000110;
filter5[7][690] = 35'b00000110101010011100111001101000000;
filter5[7][691] = 35'b11111000001011001100000111001000000;
filter5[7][692] = 35'b11111111011001000000111100100010000;
filter5[7][693] = 35'b00000100100001011000011110011000000;
filter5[7][694] = 35'b11111011011100100011001001001000000;
filter5[7][695] = 35'b00000010000111010101000010001000000;
filter5[7][696] = 35'b11111110110001010010011110010110000;
filter5[7][697] = 35'b00000011000111110010011110010000000;
filter5[7][698] = 35'b00000000101111000100100010100110000;
filter5[7][699] = 35'b11111101000100101000011111001000000;
filter5[7][700] = 35'b00000101111001100001010101001000000;
filter5[7][701] = 35'b11111011110110110110101010001000000;
filter5[7][702] = 35'b00000010101101101000010111001100000;
filter5[7][703] = 35'b00000110001100000000011000001000000;
filter5[7][704] = 35'b11111110100000100000011100110100000;
filter5[7][705] = 35'b11111111001110011001101011111000000;
filter5[7][706] = 35'b11111111100100100101010110101101000;
filter5[7][707] = 35'b11111110011001100011100000011000000;
filter5[7][708] = 35'b11111111111000000001101010010100110;
filter5[7][709] = 35'b00000000101100100100101010001000000;
filter5[7][710] = 35'b11111111000011000110111000111011000;
filter5[7][711] = 35'b00000000010000001100111100100001000;
filter5[7][712] = 35'b11111110111111001000001101100110000;
filter5[7][713] = 35'b00000000011010011001100100011100000;
filter5[7][714] = 35'b11111110101000110100001000010110000;
filter5[7][715] = 35'b11111111000001011101101100110101000;
filter5[7][716] = 35'b00000001010101000000101010010110000;
filter5[7][717] = 35'b11111101100110111001011110011100000;
filter5[7][718] = 35'b11111111101110000011001111011111100;
filter5[7][719] = 35'b11111111001000111101110010111011000;
filter5[7][720] = 35'b11111111010001101010100101000010000;
filter5[7][721] = 35'b00000000000101011001010111100001000;
filter5[7][722] = 35'b11111111110100100111000110111111000;
filter5[7][723] = 35'b11111110011100001011110001101100000;
filter5[7][724] = 35'b11111111110000101010010110110000000;
filter5[7][725] = 35'b00000000110111110010011010001101000;
filter5[7][726] = 35'b00000000101100011010110011101110000;
filter5[7][727] = 35'b00000000000111100110010111110001111;
filter5[7][728] = 35'b11111111010011100100101001011101000;
filter5[7][729] = 35'b11111110111000100000011010100110000;
filter5[7][730] = 35'b11111100111011000000001101101100000;
filter5[7][731] = 35'b00000000100010000110001101110101000;
filter5[7][732] = 35'b00000001101110101001000011000100000;
filter5[7][733] = 35'b11111110110101110001101000110100000;
filter5[7][734] = 35'b11111111010010100010101101110000000;
filter5[7][735] = 35'b11111111110000110000011101100010100;
filter5[7][736] = 35'b11111111110100101000001100010010110;
filter5[7][737] = 35'b11111111001110110110101110111110000;
filter5[7][738] = 35'b00000011000110101001011001101000000;
filter5[7][739] = 35'b11111111101010001100101000010100000;
filter5[7][740] = 35'b11111110111001010101100011010100000;
filter5[7][741] = 35'b00000001000100101001000010001100000;
filter5[7][742] = 35'b11111010111111010010000010000000000;
filter5[7][743] = 35'b11111111111000000101110011100100011;
filter5[7][744] = 35'b11111111000011011110110010111111000;
filter5[7][745] = 35'b11111111111110100011011100101001101;
filter5[7][746] = 35'b00000100110011001100111100000000000;
filter5[7][747] = 35'b11111100110111101101111100110000000;
filter5[7][748] = 35'b00000000011110011100000100011011000;
filter5[7][749] = 35'b11111111001011011110111011101011000;
filter5[7][750] = 35'b11111111010100000111010011010001000;
filter5[7][751] = 35'b11111100000110110000111111001000000;
filter5[7][752] = 35'b00000000011011001111011000000011100;
filter5[7][753] = 35'b00000000110101101101100000110101000;
filter5[7][754] = 35'b00000101000111000011100100110000000;
filter5[7][755] = 35'b11111111100101010001010101110110100;
filter5[7][756] = 35'b00000000111000010001100100110001000;
filter5[7][757] = 35'b00000100010111100100001100000000000;
filter5[7][758] = 35'b11111110101010000010101000010110000;
filter5[7][759] = 35'b11111111001101100110001101000100000;
filter5[7][760] = 35'b11111110100100011001001000001110000;
filter5[7][761] = 35'b00000000000111001101101001111110011;
filter5[7][762] = 35'b11111101011111111111101001000100000;
filter5[7][763] = 35'b11111101000100100101101100111100000;
filter5[7][764] = 35'b00000000100110111101110011111111000;
filter5[7][765] = 35'b11111110010100101111111011100000000;
filter5[7][766] = 35'b11111100010100000011111010100100000;
filter5[7][767] = 35'b11111110000010001011010001000010000;
filter5[7][768] = 35'b11111011011110111011000001100000000;
filter5[7][769] = 35'b00000010011110011001101010001000000;
filter5[7][770] = 35'b00000100010010100001101011100000000;
filter5[7][771] = 35'b00000000110110010110011010010101000;
filter5[7][772] = 35'b00000000000000111110100011100001101;
filter5[7][773] = 35'b00000000110111001011100000001100000;
filter5[7][774] = 35'b00000010110101100110011000101000000;
filter5[7][775] = 35'b00000001000001111111010011010110000;
filter5[7][776] = 35'b00000001111011000010010010101110000;
filter5[7][777] = 35'b00000001110011110111110101010110000;
filter5[7][778] = 35'b11111111100111000111101101101010100;
filter5[7][779] = 35'b00000011011111101011001110010000000;
filter5[7][780] = 35'b11111100100000111111100001001000000;
filter5[7][781] = 35'b00000010101011010100000001100000000;
filter5[7][782] = 35'b00000001100100010110001100000000000;
filter5[7][783] = 35'b00000010101110100011001011001000000;
filter5[7][784] = 35'b11111101000100101101011001010000000;
filter5[7][785] = 35'b00000011000101101001110010000100000;
filter5[7][786] = 35'b00000010000000111000011000110100000;
filter5[7][787] = 35'b11111101011001011111100101110000000;
filter5[7][788] = 35'b11111110110000111111110011111010000;
filter5[7][789] = 35'b00000011101000100000001101000100000;
filter5[7][790] = 35'b00000000101100010101001000111011000;
filter5[7][791] = 35'b00000001100000101101011100010100000;
filter5[7][792] = 35'b11111110100001101011111011111110000;
filter5[7][793] = 35'b11111111001001001010000011000001000;
filter5[7][794] = 35'b11111110000001101111011101000000000;
filter5[7][795] = 35'b00000001100110101110100010000110000;
filter5[7][796] = 35'b00000011110000000011101100110100000;
filter5[7][797] = 35'b00000000011011001010101010110000100;
filter5[7][798] = 35'b00000010001000110010110100010100000;
filter5[7][799] = 35'b11111101001111101011110010011000000;
filter5[7][800] = 35'b00000000001101010111100100000101100;
filter5[7][801] = 35'b00000001111101001000101000101110000;
filter5[7][802] = 35'b11111101100101100111111000100100000;
filter5[7][803] = 35'b00000001010100001010000001010000000;
filter5[7][804] = 35'b11111001111010010101101100001000000;
filter5[7][805] = 35'b11111111000100111001110001101111000;
filter5[7][806] = 35'b11111010101110001111100001100000000;
filter5[7][807] = 35'b11111110001000101100010111010100000;
filter5[7][808] = 35'b00000001010100010110100100101100000;
filter5[7][809] = 35'b00000110100101110011001100001000000;
filter5[7][810] = 35'b00000000101000100010010110001110000;
filter5[7][811] = 35'b11110011011001010101111101000000000;
filter5[7][812] = 35'b11111111110000110001101111110100010;
filter5[7][813] = 35'b11101110110111001000101011000000000;
filter5[7][814] = 35'b00000010010101001001111010110100000;
filter5[7][815] = 35'b00000101011001001111010010111000000;
filter5[7][816] = 35'b00000000010100100011001111100010100;
filter5[7][817] = 35'b11111111110011111111000000111011100;
filter5[7][818] = 35'b00001010100100110010101010110000000;
filter5[7][819] = 35'b11111010110110110101100111110000000;
filter5[7][820] = 35'b11110110111111100100000010000000000;
filter5[7][821] = 35'b00001000000111101010110000000000000;
filter5[7][822] = 35'b00000000100010101010011110001111000;
filter5[7][823] = 35'b11111111111110011110010110111010111;
filter5[7][824] = 35'b00000000111011001010011101100111000;
filter5[7][825] = 35'b00000000001110011010001101000100010;
filter5[7][826] = 35'b11111110010001000011101101011100000;
filter5[7][827] = 35'b11111011011010110110010110100000000;
filter5[7][828] = 35'b11111110100110000011010110100110000;
filter5[7][829] = 35'b00000001011101100011110110011110000;
filter5[7][830] = 35'b11111110110001110011101001101000000;
filter5[7][831] = 35'b00000001000110101011100000011010000;
filter5[7][832] = 35'b11111110101100001010110110101000000;
filter5[7][833] = 35'b11111111011100101011111011100010000;
filter5[7][834] = 35'b11111101111110011101110111001000000;
filter5[7][835] = 35'b11111110001100001110001100011000000;
filter5[7][836] = 35'b11111111001001000101101100011010000;
filter5[7][837] = 35'b00000000001010111000010011111001000;
filter5[7][838] = 35'b11111110101110000010111000010100000;
filter5[7][839] = 35'b00000000000110001101010010110001100;
filter5[7][840] = 35'b11111111100011001100111010111100100;
filter5[7][841] = 35'b11111110100100000101000000011100000;
filter5[7][842] = 35'b11111111010100111111110111100110000;
filter5[7][843] = 35'b11111110011010101100100011001110000;
filter5[7][844] = 35'b11111111111110100110001101100101101;
filter5[7][845] = 35'b11111111101001101101111001110001000;
filter5[7][846] = 35'b11111111100110010101111111110011000;
filter5[7][847] = 35'b00000000010010010010011010101000000;
filter5[7][848] = 35'b11111111011001110100110100110010000;
filter5[7][849] = 35'b00000000011001110001010101011011100;
filter5[7][850] = 35'b11111111110001100100100111101010100;
filter5[7][851] = 35'b00000000101000010001001000011001000;
filter5[7][852] = 35'b00000001001011100001001100110000000;
filter5[7][853] = 35'b11111101101101101001001011110100000;
filter5[7][854] = 35'b11111110100010000101010000010100000;
filter5[7][855] = 35'b11111111011111110100100001101011000;
filter5[7][856] = 35'b11111111000011100010000000010111000;
filter5[7][857] = 35'b11111110110111110101011000110010000;
filter5[7][858] = 35'b00000000100110001011000100111000000;
filter5[7][859] = 35'b11111011010001111101001100101000000;
filter5[7][860] = 35'b11111101011010110010011000010000000;
filter5[7][861] = 35'b11111110110110110011101101111000000;
filter5[7][862] = 35'b00000001010111100110111100111010000;
filter5[7][863] = 35'b11111111111010111101010110000010000;
filter5[7][864] = 35'b00000001000011101000101011000110000;
filter5[7][865] = 35'b11111110111110101100001001111000000;
filter5[7][866] = 35'b00000001101101111010100000111100000;
filter5[7][867] = 35'b11111111100011110111101101000110100;
filter5[7][868] = 35'b00000000011011000111101001101000100;
filter5[7][869] = 35'b00000010011100000101010010110000000;
filter5[7][870] = 35'b11111101011111000011110110000100000;
filter5[7][871] = 35'b11111111110111110111001111000111100;
filter5[7][872] = 35'b11111111101110111111000111101100000;
filter5[7][873] = 35'b11111100011011001000011101111000000;
filter5[7][874] = 35'b11111011101111100001010110000000000;
filter5[7][875] = 35'b11111101000010000001010111011000000;
filter5[7][876] = 35'b00000010011100111100000101111100000;
filter5[7][877] = 35'b00000100110001100001011100000000000;
filter5[7][878] = 35'b00000001111100010101100001100110000;
filter5[7][879] = 35'b11111011001001110110101100010000000;
filter5[7][880] = 35'b00000001100110101101110101100000000;
filter5[7][881] = 35'b00000010111001110001111011111100000;
filter5[7][882] = 35'b00000011011010001101001000101000000;
filter5[7][883] = 35'b00000001010111010101110110111100000;
filter5[7][884] = 35'b11111111101101111110010111101011100;
filter5[7][885] = 35'b00000000110110100010011010100100000;
filter5[7][886] = 35'b11110110011000111100111110000000000;
filter5[7][887] = 35'b00000000011011100000101111010110100;
filter5[7][888] = 35'b00000001000000001100110010111010000;
filter5[7][889] = 35'b11111101111110001010000000111100000;
filter5[7][890] = 35'b00000000110101111111011011110111000;
filter5[7][891] = 35'b00000001101110110000010010001010000;
filter5[7][892] = 35'b11111110010011011000111111100000000;
filter5[7][893] = 35'b11111110000001011010110000011000000;
filter5[7][894] = 35'b11111101011011011101111100000000000;
filter5[7][895] = 35'b11111110110111101001011110111110000;
filter5[7][896] = 35'b00000010001000100100111110010100000;
filter5[7][897] = 35'b11111010010001111101110111010000000;
filter5[7][898] = 35'b00001000000110000101111000010000000;
filter5[7][899] = 35'b00000010010100001100100111010000000;
filter5[7][900] = 35'b00001001101101000001011000100000000;
filter5[7][901] = 35'b11111011100001011110000011110000000;
filter5[7][902] = 35'b00000000001110000101101010101100110;
filter5[7][903] = 35'b00000101100110101010111000101000000;
filter5[7][904] = 35'b11111100010001000110011010100100000;
filter5[7][905] = 35'b11111101100111110010101000101000000;
filter5[7][906] = 35'b00000011111110101010010001111000000;
filter5[7][907] = 35'b11111101001100101101011111110100000;
filter5[7][908] = 35'b11110101100110110101000000100000000;
filter5[7][909] = 35'b11111100100000101011010110100000000;
filter5[7][910] = 35'b00000011010100010100101110011100000;
filter5[7][911] = 35'b00000011101111000110100010101100000;
filter5[7][912] = 35'b11111100100101001010011100111000000;
filter5[7][913] = 35'b11110110011010110001010100010000000;
filter5[7][914] = 35'b11111100110000000010111101101000000;
filter5[7][915] = 35'b11111100111011010110010001110000000;
filter5[7][916] = 35'b00000001110100000110010110000010000;
filter5[7][917] = 35'b11101101111110100001111100000000000;
filter5[7][918] = 35'b11111010110011100101110011100000000;
filter5[7][919] = 35'b00000110011011010011101100011000000;
filter5[7][920] = 35'b11110000110010101100011101100000000;
filter5[7][921] = 35'b11110100011101011101100001010000000;
filter5[7][922] = 35'b11110111101010001011100000110000000;
filter5[7][923] = 35'b00000000111011100101001111111111000;
filter5[7][924] = 35'b11111011010111001001010010001000000;
filter5[7][925] = 35'b11111010111110001001001010011000000;
filter5[7][926] = 35'b11101110111000101101101101100000000;
filter5[7][927] = 35'b11111111110111000010101010010111110;
filter5[7][928] = 35'b00000001010010100000010111010010000;
filter5[7][929] = 35'b11111010110111111010010110011000000;
filter5[7][930] = 35'b00000011100100110101101101011100000;
filter5[7][931] = 35'b00000011100101101010101110011100000;
filter5[7][932] = 35'b11111110111011101000100100111010000;
filter5[7][933] = 35'b11111110111001001010110011010000000;
filter5[7][934] = 35'b11110010111011000101101101110000000;
filter5[7][935] = 35'b11111000111110000000110000010000000;
filter5[7][936] = 35'b11111101101101100010000101001100000;
filter5[7][937] = 35'b11111101000111001101100010000000000;
filter5[7][938] = 35'b00000001100001010000011110001000000;
filter5[7][939] = 35'b11111011100010001101011100011000000;
filter5[7][940] = 35'b11111110010100111011000001000000000;
filter5[7][941] = 35'b00000110100001011010001101001000000;
filter5[7][942] = 35'b00000010011100010010101111001000000;
filter5[7][943] = 35'b11110101010010110101110000010000000;
filter5[7][944] = 35'b00000010000101110001111100000000000;
filter5[7][945] = 35'b00000100111001111101000001111000000;
filter5[7][946] = 35'b11111100011011010011101101110000000;
filter5[7][947] = 35'b11111110010100110100111001111110000;
filter5[7][948] = 35'b00000100110011001011101110110000000;
filter5[7][949] = 35'b11111110000010010100101110010000000;
filter5[7][950] = 35'b11110001111011011010001000000000000;
filter5[7][951] = 35'b11111100000000010110011001010000000;
filter5[7][952] = 35'b11111111111011000011011010010000010;
filter5[7][953] = 35'b11100110011111000011110001100000000;
filter5[7][954] = 35'b11111010000000001001101000101000000;
filter5[7][955] = 35'b00000000000010011110111001110101000;
filter5[7][956] = 35'b00000100111111111101111111110000000;
filter5[7][957] = 35'b00000010001111000101101111000000000;
filter5[7][958] = 35'b11101111011011100101011001100000000;
filter5[7][959] = 35'b11111011111011011011110010010000000;
filter5[7][960] = 35'b11111111010000011010001000111001000;
filter5[7][961] = 35'b00000001010000111101101101100010000;
filter5[7][962] = 35'b11111010110000111011010001000000000;
filter5[7][963] = 35'b00001010000100111110000101100000000;
filter5[7][964] = 35'b00001000101000001001111100010000000;
filter5[7][965] = 35'b00001000001000011101101110100000000;
filter5[7][966] = 35'b00000001000001100111111001011110000;
filter5[7][967] = 35'b00000101001000000111110110101000000;
filter5[7][968] = 35'b00000100101100110011001000010000000;
filter5[7][969] = 35'b00000001110110011100100101110100000;
filter5[7][970] = 35'b11111111000011101000110101110001000;
filter5[7][971] = 35'b00000000111111101011110100001110000;
filter5[7][972] = 35'b00000001111001011011011100111010000;
filter5[7][973] = 35'b00000010111011010010111110111000000;
filter5[7][974] = 35'b00000011001011100101000010101000000;
filter5[7][975] = 35'b00000001101110111000001111001010000;
filter5[7][976] = 35'b11111110010001110001111001000000000;
filter5[7][977] = 35'b11111101001011000111001000001000000;
filter5[7][978] = 35'b11110011110001111111010001000000000;
filter5[7][979] = 35'b00000010111011001000100000111100000;
filter5[7][980] = 35'b11111110011101010011010110010100000;
filter5[7][981] = 35'b00000000110110010011110010000110000;
filter5[7][982] = 35'b11111001010110011101100101100000000;
filter5[7][983] = 35'b11111000011011110111100111001000000;
filter5[7][984] = 35'b11111100111110101011011010010000000;
filter5[7][985] = 35'b00000010000110001010011100011100000;
filter5[7][986] = 35'b11111001111000100100001010011000000;
filter5[7][987] = 35'b11111100100110000000011010101000000;
filter5[7][988] = 35'b11111111001010001010001100110111000;
filter5[7][989] = 35'b11111011101010011010010111110000000;
filter5[7][990] = 35'b00000000110001110111001001110110000;
filter5[7][991] = 35'b11111101010001001010011000011100000;
filter5[7][992] = 35'b11111010100000111111100000010000000;
filter5[7][993] = 35'b00000000100100000100011010000000000;
filter5[7][994] = 35'b00000110011100011001100100110000000;
filter5[7][995] = 35'b00000001100010011001101001010110000;
filter5[7][996] = 35'b00000000110110101001010110010111000;
filter5[7][997] = 35'b11111110000000110110101110110010000;
filter5[7][998] = 35'b00000100001101111111010111111000000;
filter5[7][999] = 35'b11110001000000001001010101010000000;
filter5[7][1000] = 35'b11111010110101010000111110000000000;
filter5[7][1001] = 35'b11111100100011100110000101000000000;
filter5[7][1002] = 35'b00000001010110001101001010000100000;
filter5[7][1003] = 35'b11111110110011000100010010111010000;
filter5[7][1004] = 35'b00000001100001111100110000100000000;
filter5[7][1005] = 35'b00000000101111001111000000100001000;
filter5[7][1006] = 35'b00000001000111000011101101100000000;
filter5[7][1007] = 35'b00000001010001101010000000110000000;
filter5[7][1008] = 35'b00000000111001110111010110101000000;
filter5[7][1009] = 35'b00000010100101001000011101110100000;
filter5[7][1010] = 35'b00001100101111110001111101110000000;
filter5[7][1011] = 35'b11111100111000101111000111001000000;
filter5[7][1012] = 35'b00000011011000110101110100000100000;
filter5[7][1013] = 35'b11111101011011101011001110110100000;
filter5[7][1014] = 35'b00000011100110110001100110000100000;
filter5[7][1015] = 35'b11111100100100011001101001011100000;
filter5[7][1016] = 35'b11111100110111111000100010101000000;
filter5[7][1017] = 35'b11111110000110001001111001101110000;
filter5[7][1018] = 35'b11111001110011010101101101010000000;
filter5[7][1019] = 35'b11111100100111111001001111111100000;
filter5[7][1020] = 35'b00000101110101110000010111100000000;
filter5[7][1021] = 35'b11110101111000001010001010110000000;
filter5[7][1022] = 35'b11110111001101011100110010000000000;
filter5[7][1023] = 35'b11111111011000001101110111010010000;
filter5[8][0] = 35'b00000000110001011001110110110000000;
filter5[8][1] = 35'b00000011011101010101001011000100000;
filter5[8][2] = 35'b11111111011011010010011101010100000;
filter5[8][3] = 35'b11111100010000110000011110111000000;
filter5[8][4] = 35'b11111101001000010111101100101100000;
filter5[8][5] = 35'b11111101010101110000000011101100000;
filter5[8][6] = 35'b11111111101100000011000100101010100;
filter5[8][7] = 35'b00000000101011010100110010010010000;
filter5[8][8] = 35'b00000010110010101001110001001100000;
filter5[8][9] = 35'b11111011100001001100001101110000000;
filter5[8][10] = 35'b11111111111000111001100100100101101;
filter5[8][11] = 35'b00000011100110110111000110110100000;
filter5[8][12] = 35'b11111011101101000101011101101000000;
filter5[8][13] = 35'b00000100011100000001010101101000000;
filter5[8][14] = 35'b00000111011000111010001011100000000;
filter5[8][15] = 35'b00000111100010110000001011001000000;
filter5[8][16] = 35'b11111111011000100001000001110011000;
filter5[8][17] = 35'b11111111010110111100011110001101000;
filter5[8][18] = 35'b11111001100000100111001111111000000;
filter5[8][19] = 35'b00000010001011100110100010000000000;
filter5[8][20] = 35'b00000001101100000000111011111010000;
filter5[8][21] = 35'b11111101001101110101101100111000000;
filter5[8][22] = 35'b00000111001001011010110011001000000;
filter5[8][23] = 35'b00000100100100111001111111011000000;
filter5[8][24] = 35'b00000011111011010110000010111100000;
filter5[8][25] = 35'b00000000101001100111111001110110000;
filter5[8][26] = 35'b11111111110001011011101000010000000;
filter5[8][27] = 35'b00000001100101111011011010001000000;
filter5[8][28] = 35'b11111111100010100111000110111011100;
filter5[8][29] = 35'b11111011001100100001111001110000000;
filter5[8][30] = 35'b00000010001111000111000010101100000;
filter5[8][31] = 35'b11111100100101001111000101111100000;
filter5[8][32] = 35'b11111111001100111001001111111111000;
filter5[8][33] = 35'b00000001001110000101110011110010000;
filter5[8][34] = 35'b00000010010100001000101111011000000;
filter5[8][35] = 35'b11111100010000011100101100101000000;
filter5[8][36] = 35'b00000001100110010111010100111010000;
filter5[8][37] = 35'b00000010010001011001001001010100000;
filter5[8][38] = 35'b11101111100011010010110010100000000;
filter5[8][39] = 35'b11111000101101100101110001100000000;
filter5[8][40] = 35'b00000010000011111001001010111100000;
filter5[8][41] = 35'b11111111101100100100110111000010100;
filter5[8][42] = 35'b11111110100100010001010000111110000;
filter5[8][43] = 35'b00000100111000010111001011001000000;
filter5[8][44] = 35'b00000011011101000101011101010100000;
filter5[8][45] = 35'b11111011011000111110101101000000000;
filter5[8][46] = 35'b11110110011110100111000111000000000;
filter5[8][47] = 35'b00000001110000111101000011110110000;
filter5[8][48] = 35'b00000000111010101110110100111110000;
filter5[8][49] = 35'b11111110100010011101110001011100000;
filter5[8][50] = 35'b00000011111101001110011111111100000;
filter5[8][51] = 35'b11111100100101010111010000011000000;
filter5[8][52] = 35'b11111110000110111101011100000010000;
filter5[8][53] = 35'b11110011110000001100101100100000000;
filter5[8][54] = 35'b11111110101101011010010110100000000;
filter5[8][55] = 35'b11111101001101010111001010010000000;
filter5[8][56] = 35'b11111111001000001011001101011110000;
filter5[8][57] = 35'b11111110110100101011000101001100000;
filter5[8][58] = 35'b11111100101011011011000111100000000;
filter5[8][59] = 35'b00000000110111101101000000101000000;
filter5[8][60] = 35'b00000100011101111000011011110000000;
filter5[8][61] = 35'b11111010100010100001011111111000000;
filter5[8][62] = 35'b00000001010000000101100011001100000;
filter5[8][63] = 35'b00000001010100001110001101011100000;
filter5[8][64] = 35'b00000001010001101011101011100010000;
filter5[8][65] = 35'b11111101001001000010000001011100000;
filter5[8][66] = 35'b00000001101001000110010100010100000;
filter5[8][67] = 35'b11111001011011011110011010010000000;
filter5[8][68] = 35'b11111111101001101000000110011001100;
filter5[8][69] = 35'b11111011111101101111000100010000000;
filter5[8][70] = 35'b00000000111011101010010010000001000;
filter5[8][71] = 35'b00000001010000110010110011110000000;
filter5[8][72] = 35'b00000001010010111001001101110100000;
filter5[8][73] = 35'b11111111110000010111100111000101010;
filter5[8][74] = 35'b11111100110101100111111111100000000;
filter5[8][75] = 35'b00000001111011110101011100111010000;
filter5[8][76] = 35'b11111001011100011100110110000000000;
filter5[8][77] = 35'b11111101100001011110011100001100000;
filter5[8][78] = 35'b00000100010110001001001101110000000;
filter5[8][79] = 35'b00000001100110011001011100010000000;
filter5[8][80] = 35'b11111111011101011100110101001010000;
filter5[8][81] = 35'b11111111111101001010010101011101101;
filter5[8][82] = 35'b11111010000110100110111000110000000;
filter5[8][83] = 35'b00000001011000101110000010111000000;
filter5[8][84] = 35'b00000000111111100011101001001111000;
filter5[8][85] = 35'b00000000111011000000101010010000000;
filter5[8][86] = 35'b11111100111011010001001010111100000;
filter5[8][87] = 35'b00000001100101000000101100010110000;
filter5[8][88] = 35'b00000001000100100011011000011000000;
filter5[8][89] = 35'b11111101100001100000100110010100000;
filter5[8][90] = 35'b11111110010010100111000011010000000;
filter5[8][91] = 35'b00000000110010111110101110010100000;
filter5[8][92] = 35'b11111110110011100000111010011010000;
filter5[8][93] = 35'b11111100011101011111011001100100000;
filter5[8][94] = 35'b11111110111100110101010010101110000;
filter5[8][95] = 35'b00000001000111010111100101110000000;
filter5[8][96] = 35'b11111011010010111010101111001000000;
filter5[8][97] = 35'b00000000110001001101010111101110000;
filter5[8][98] = 35'b00000100010001111100010000100000000;
filter5[8][99] = 35'b11111111111111011111111010001000011;
filter5[8][100] = 35'b00000000111010010100100001100111000;
filter5[8][101] = 35'b11111100111001011110000110111100000;
filter5[8][102] = 35'b11111101101001111101110011101000000;
filter5[8][103] = 35'b11111101100110011101100111101100000;
filter5[8][104] = 35'b11111111100011000001101111101101100;
filter5[8][105] = 35'b11111111101010000100111010010110000;
filter5[8][106] = 35'b11111101111110011110110110111100000;
filter5[8][107] = 35'b00000001010111000111101101011110000;
filter5[8][108] = 35'b00000000011011010010000010000011000;
filter5[8][109] = 35'b11111111010111111001101001101000000;
filter5[8][110] = 35'b11111011111110101110011010011000000;
filter5[8][111] = 35'b00000010010111100110111011011100000;
filter5[8][112] = 35'b11111101011011010001110110100100000;
filter5[8][113] = 35'b00000001111010111110110000011110000;
filter5[8][114] = 35'b00000001011101110000000111010110000;
filter5[8][115] = 35'b11111110110011000011010110101000000;
filter5[8][116] = 35'b00000000101000001001111010010101000;
filter5[8][117] = 35'b00000100000011100000001010001000000;
filter5[8][118] = 35'b00000000000011000001010110000110110;
filter5[8][119] = 35'b11111100111011010010000100101000000;
filter5[8][120] = 35'b00000010111111010011111101100100000;
filter5[8][121] = 35'b11111001001111101001000010100000000;
filter5[8][122] = 35'b11111010000101011000010110100000000;
filter5[8][123] = 35'b00000010000011101111000110001100000;
filter5[8][124] = 35'b00000000100001000001101000000101000;
filter5[8][125] = 35'b00000101110110111011110010100000000;
filter5[8][126] = 35'b11110101111101001011001010010000000;
filter5[8][127] = 35'b11111101111111001110011111001100000;
filter5[8][128] = 35'b11110101001010110111111000100000000;
filter5[8][129] = 35'b11101101011100010011110111000000000;
filter5[8][130] = 35'b00000000100001001000001101101001000;
filter5[8][131] = 35'b11101111100001100110011000100000000;
filter5[8][132] = 35'b11111111001100110101001010101111000;
filter5[8][133] = 35'b11111000110101111000101110010000000;
filter5[8][134] = 35'b11111010111101111011011100011000000;
filter5[8][135] = 35'b00000010110110000001101101110000000;
filter5[8][136] = 35'b00000000010101111011010001001101000;
filter5[8][137] = 35'b11111000110100100111000101001000000;
filter5[8][138] = 35'b11110001111010111000100000010000000;
filter5[8][139] = 35'b11110101001010101101011001010000000;
filter5[8][140] = 35'b11101000010101001110101111100000000;
filter5[8][141] = 35'b11101110101110110110111010100000000;
filter5[8][142] = 35'b00000011000000111011010010111100000;
filter5[8][143] = 35'b11111001100111000010010110010000000;
filter5[8][144] = 35'b11110111110111001100111111100000000;
filter5[8][145] = 35'b11110001001111011111111110110000000;
filter5[8][146] = 35'b11111000001100111000001011110000000;
filter5[8][147] = 35'b11111111101001000000000111101111100;
filter5[8][148] = 35'b00000010011010011111111000011000000;
filter5[8][149] = 35'b11111100100000100101000001101100000;
filter5[8][150] = 35'b11100110000001011110000010000000000;
filter5[8][151] = 35'b11111100000101011100011011111100000;
filter5[8][152] = 35'b11111011100001010100110111110000000;
filter5[8][153] = 35'b11111000111011001011001110110000000;
filter5[8][154] = 35'b11111110011011100000000000001010000;
filter5[8][155] = 35'b11111110111100101000011011110010000;
filter5[8][156] = 35'b11111010000110111010000010010000000;
filter5[8][157] = 35'b00000110001001010001000000010000000;
filter5[8][158] = 35'b00000001011111101010001011100010000;
filter5[8][159] = 35'b11111111100011011000011001110000100;
filter5[8][160] = 35'b11110111011001100011011000010000000;
filter5[8][161] = 35'b00001000010111100010010101010000000;
filter5[8][162] = 35'b11111110111011011101111010110100000;
filter5[8][163] = 35'b00000000101001111100010000101111000;
filter5[8][164] = 35'b11111000111000001011011010001000000;
filter5[8][165] = 35'b00000001011000001000100101001010000;
filter5[8][166] = 35'b11111101001100111110000101111100000;
filter5[8][167] = 35'b11111100110101100111001010011100000;
filter5[8][168] = 35'b11110110101011100100110011100000000;
filter5[8][169] = 35'b11111110111001000100110010000110000;
filter5[8][170] = 35'b11111010110001110001010110111000000;
filter5[8][171] = 35'b00000000010011100001110000010101100;
filter5[8][172] = 35'b00000000111010100000000000011000000;
filter5[8][173] = 35'b00000101100011110110111100010000000;
filter5[8][174] = 35'b00000000000111101011101011110101111;
filter5[8][175] = 35'b11111100110110101100000101101100000;
filter5[8][176] = 35'b00000101000110000001100010111000000;
filter5[8][177] = 35'b00000001101101111110111101000010000;
filter5[8][178] = 35'b11111001001110010101011000010000000;
filter5[8][179] = 35'b11111000010100000100101001011000000;
filter5[8][180] = 35'b00000010100011010010100110111100000;
filter5[8][181] = 35'b00001101010001100000000010000000000;
filter5[8][182] = 35'b11110001001100010101101001100000000;
filter5[8][183] = 35'b00000011110010101001001110000100000;
filter5[8][184] = 35'b11111010011000111011000010101000000;
filter5[8][185] = 35'b00000001001101101100110100000010000;
filter5[8][186] = 35'b11101000011111110011110001000000000;
filter5[8][187] = 35'b11111010101000101110000101110000000;
filter5[8][188] = 35'b00001011101110100100001111100000000;
filter5[8][189] = 35'b11111101110001100101110101110000000;
filter5[8][190] = 35'b11110101010010111001110111110000000;
filter5[8][191] = 35'b11101100000111010001010000000000000;
filter5[8][192] = 35'b11111000110010001100001111101000000;
filter5[8][193] = 35'b11111111001100010011111100001010000;
filter5[8][194] = 35'b11110100111010101110101001000000000;
filter5[8][195] = 35'b00000001001001100111100001111010000;
filter5[8][196] = 35'b11110100000111011100101010010000000;
filter5[8][197] = 35'b11111000100000001011111001111000000;
filter5[8][198] = 35'b11111100010111100111011101000100000;
filter5[8][199] = 35'b11111111011011001011100000001101000;
filter5[8][200] = 35'b11111000111110000100000001110000000;
filter5[8][201] = 35'b11111000110110011110111011000000000;
filter5[8][202] = 35'b00000111001011111010011011111000000;
filter5[8][203] = 35'b11111100101000000011110000101000000;
filter5[8][204] = 35'b11111101011100101101001011011100000;
filter5[8][205] = 35'b11111110110100110010000000111110000;
filter5[8][206] = 35'b00000001010001110000001011010010000;
filter5[8][207] = 35'b11111101011011100011011101101000000;
filter5[8][208] = 35'b11111011111011010000101010000000000;
filter5[8][209] = 35'b00000110000110000000110000001000000;
filter5[8][210] = 35'b11110111111010111110110111110000000;
filter5[8][211] = 35'b11101011000111110010001011000000000;
filter5[8][212] = 35'b11111110011111011100111111011100000;
filter5[8][213] = 35'b11111100101001110001111110011000000;
filter5[8][214] = 35'b00000011011001011100101111100000000;
filter5[8][215] = 35'b11111000110001100000000110100000000;
filter5[8][216] = 35'b11111110110011100011111101000110000;
filter5[8][217] = 35'b11111001110011011101010110110000000;
filter5[8][218] = 35'b11110101111100101000111000010000000;
filter5[8][219] = 35'b11111111110010101100111001101100010;
filter5[8][220] = 35'b00000010100101001111011011011100000;
filter5[8][221] = 35'b00000010111001110100011100010100000;
filter5[8][222] = 35'b11111101001001100100110000110100000;
filter5[8][223] = 35'b00000100001010110010010101001000000;
filter5[8][224] = 35'b00010000111101001001010110000000000;
filter5[8][225] = 35'b11111101110011101101100111001000000;
filter5[8][226] = 35'b11111001010011110000001111010000000;
filter5[8][227] = 35'b00000100110111111011111001101000000;
filter5[8][228] = 35'b11111010010011111001000000010000000;
filter5[8][229] = 35'b00000100000110110110001010000000000;
filter5[8][230] = 35'b11111010000100011110111000110000000;
filter5[8][231] = 35'b11111001110000011110100010111000000;
filter5[8][232] = 35'b11110110101110010011010100000000000;
filter5[8][233] = 35'b00000100011010111101001110100000000;
filter5[8][234] = 35'b11111101110001011000101110011100000;
filter5[8][235] = 35'b11111100010011101100111100100000000;
filter5[8][236] = 35'b00000000010000010111011110011100100;
filter5[8][237] = 35'b00000000101010110101110100110101000;
filter5[8][238] = 35'b11111111010010000101100110111110000;
filter5[8][239] = 35'b11111011111011011001110100101000000;
filter5[8][240] = 35'b11101101000001101000011100100000000;
filter5[8][241] = 35'b11111101011110000011000001001100000;
filter5[8][242] = 35'b00000110101001001011111111000000000;
filter5[8][243] = 35'b11111111101011100101100101100100000;
filter5[8][244] = 35'b11111101101101110100100010101100000;
filter5[8][245] = 35'b00000010100110100101111010010100000;
filter5[8][246] = 35'b11111111101101001000011000011111000;
filter5[8][247] = 35'b11111010010001110111111110011000000;
filter5[8][248] = 35'b11111101110001111001000111010000000;
filter5[8][249] = 35'b11111010110111100100110100110000000;
filter5[8][250] = 35'b00001000111011010010000111100000000;
filter5[8][251] = 35'b11111010101001100011110001101000000;
filter5[8][252] = 35'b00000001010001110101010111111100000;
filter5[8][253] = 35'b00000101000011010011000011100000000;
filter5[8][254] = 35'b11111011001110011000101100101000000;
filter5[8][255] = 35'b11111000101001011101110011100000000;
filter5[8][256] = 35'b11111101011000100011100010011100000;
filter5[8][257] = 35'b11111111011111100100100100000101000;
filter5[8][258] = 35'b11111111000011110011001110000000000;
filter5[8][259] = 35'b11111100110100011110001010011000000;
filter5[8][260] = 35'b11111111011001111101011010010111000;
filter5[8][261] = 35'b11111111100101111111011101100010000;
filter5[8][262] = 35'b11111011110011001010110011110000000;
filter5[8][263] = 35'b11111111001110100100001100000000000;
filter5[8][264] = 35'b11111101011101010010101111111100000;
filter5[8][265] = 35'b11111111000011100111110101110100000;
filter5[8][266] = 35'b11111011101011000010000101000000000;
filter5[8][267] = 35'b11111101100110101010010101101000000;
filter5[8][268] = 35'b11111110110110100011111100001000000;
filter5[8][269] = 35'b00000010101111111100000111000000000;
filter5[8][270] = 35'b11111101111010101010001011011000000;
filter5[8][271] = 35'b11111100011000101011001010001100000;
filter5[8][272] = 35'b11111100101000010101110010101000000;
filter5[8][273] = 35'b11111010101010011010010110001000000;
filter5[8][274] = 35'b11110011100001100011100100100000000;
filter5[8][275] = 35'b11111011011011011000111100100000000;
filter5[8][276] = 35'b11111011111000000101010001001000000;
filter5[8][277] = 35'b11110010111011001001001001010000000;
filter5[8][278] = 35'b11111010000110000101110011101000000;
filter5[8][279] = 35'b11111000101001010001000001110000000;
filter5[8][280] = 35'b11110010011000001100110000000000000;
filter5[8][281] = 35'b11110111100000011100010010000000000;
filter5[8][282] = 35'b00000101011001110101010111110000000;
filter5[8][283] = 35'b11111011111001111101101101011000000;
filter5[8][284] = 35'b00000011000100001100011011001100000;
filter5[8][285] = 35'b11111100011011000011010111100000000;
filter5[8][286] = 35'b00000111110011001000010001010000000;
filter5[8][287] = 35'b11110110111110000000010101110000000;
filter5[8][288] = 35'b00001011100111001000010111110000000;
filter5[8][289] = 35'b11111101100001000010100001110000000;
filter5[8][290] = 35'b11111001011111101011101101101000000;
filter5[8][291] = 35'b00000000000010010111010000011001011;
filter5[8][292] = 35'b11111010111110011001110001000000000;
filter5[8][293] = 35'b00000100001010111011000001100000000;
filter5[8][294] = 35'b00000010100111110000000000100000000;
filter5[8][295] = 35'b11111000100011011001110101100000000;
filter5[8][296] = 35'b11110111001010010010111010000000000;
filter5[8][297] = 35'b00000100001101110111100000111000000;
filter5[8][298] = 35'b11111010111111011110000000111000000;
filter5[8][299] = 35'b00000001001000001100001001000100000;
filter5[8][300] = 35'b00000010001110100001110101001100000;
filter5[8][301] = 35'b11111111011001010100101001001011000;
filter5[8][302] = 35'b00000000001110100110011111011101010;
filter5[8][303] = 35'b11110101101100110010000101000000000;
filter5[8][304] = 35'b11111000010100100111010010000000000;
filter5[8][305] = 35'b11111100111001011101011000000100000;
filter5[8][306] = 35'b00000010001000000110010111011000000;
filter5[8][307] = 35'b00000000011010010001101011001110000;
filter5[8][308] = 35'b11111111000000000010001110000111000;
filter5[8][309] = 35'b11111110011000111001111110111010000;
filter5[8][310] = 35'b00000011001101111111100110100000000;
filter5[8][311] = 35'b11111010111010110000101001101000000;
filter5[8][312] = 35'b11111011010100101111010011000000000;
filter5[8][313] = 35'b11110110110111001010010010010000000;
filter5[8][314] = 35'b00000000101111100100110000100001000;
filter5[8][315] = 35'b00000100011110001001110101011000000;
filter5[8][316] = 35'b11111111110111001110011011111000000;
filter5[8][317] = 35'b00000011101101100000110101111100000;
filter5[8][318] = 35'b11111111000110001101100000110010000;
filter5[8][319] = 35'b11111010011011001011011011000000000;
filter5[8][320] = 35'b11111011110001001100110011111000000;
filter5[8][321] = 35'b00000001101010010100100001010000000;
filter5[8][322] = 35'b00000001100111000001111010001100000;
filter5[8][323] = 35'b00000001111000001010001100010100000;
filter5[8][324] = 35'b11111100011010101110111110101000000;
filter5[8][325] = 35'b00001000001011101011011100010000000;
filter5[8][326] = 35'b00000011101010100111001101011000000;
filter5[8][327] = 35'b00001011100001011111001001010000000;
filter5[8][328] = 35'b11111111111100100010110100010001010;
filter5[8][329] = 35'b11111011000001010001101110100000000;
filter5[8][330] = 35'b00000011000010100100110100000100000;
filter5[8][331] = 35'b00000000000111010100101001011010101;
filter5[8][332] = 35'b11111111100000001001110010110111000;
filter5[8][333] = 35'b00000000001100010111100110001011010;
filter5[8][334] = 35'b00001000010001101000000101010000000;
filter5[8][335] = 35'b00000001100011010001011000011100000;
filter5[8][336] = 35'b11111110000110111101001001001000000;
filter5[8][337] = 35'b11111101011001101100011000011000000;
filter5[8][338] = 35'b11111010001111001010010000011000000;
filter5[8][339] = 35'b00000000011011110001010000001011100;
filter5[8][340] = 35'b00000000110111111001100110011000000;
filter5[8][341] = 35'b11111101110010100111111000111000000;
filter5[8][342] = 35'b00000100010100011011010001010000000;
filter5[8][343] = 35'b00000100011000100100011011101000000;
filter5[8][344] = 35'b00000100110110000001001011001000000;
filter5[8][345] = 35'b11111111110000101110110100111011100;
filter5[8][346] = 35'b00000011110011011110101101011000000;
filter5[8][347] = 35'b00000001001100110011000000000010000;
filter5[8][348] = 35'b11111111010011100100110000101111000;
filter5[8][349] = 35'b00000001011100001000010110000000000;
filter5[8][350] = 35'b00000000001000011100111111001111010;
filter5[8][351] = 35'b11111011111110110110111010001000000;
filter5[8][352] = 35'b11111111100100110111001100001100100;
filter5[8][353] = 35'b00000001001010101011010001000110000;
filter5[8][354] = 35'b11111110000010101101111001000010000;
filter5[8][355] = 35'b11111111010000111110001100010001000;
filter5[8][356] = 35'b00000000011111001110100111011111100;
filter5[8][357] = 35'b11111111011011101111110100011101000;
filter5[8][358] = 35'b11111010010101110010011111100000000;
filter5[8][359] = 35'b11111111001010001110111101100100000;
filter5[8][360] = 35'b11111111010011110011011010111000000;
filter5[8][361] = 35'b00000001011001011111101000100100000;
filter5[8][362] = 35'b00000001100100100001011101100010000;
filter5[8][363] = 35'b00000010010110010110110110100100000;
filter5[8][364] = 35'b11111111101011001001010101110001100;
filter5[8][365] = 35'b11111111001000110110101110100101000;
filter5[8][366] = 35'b11111110110010010001011001000100000;
filter5[8][367] = 35'b11111110010111000100011011101100000;
filter5[8][368] = 35'b00000010000110110110110010110000000;
filter5[8][369] = 35'b11111101001000000000100100111000000;
filter5[8][370] = 35'b00000001100010110110000100011000000;
filter5[8][371] = 35'b00000000111110111100010101100111000;
filter5[8][372] = 35'b11111110100111011011011000101000000;
filter5[8][373] = 35'b11111111101101000010010010011101100;
filter5[8][374] = 35'b00000001100011110100111001101100000;
filter5[8][375] = 35'b11111101011010110000000001011100000;
filter5[8][376] = 35'b11111101001001011110011111101000000;
filter5[8][377] = 35'b11111010010110100011100010011000000;
filter5[8][378] = 35'b11111100000011110101000000101000000;
filter5[8][379] = 35'b11111100111100110111100110101000000;
filter5[8][380] = 35'b11111111011110100110101100100011000;
filter5[8][381] = 35'b00000011110111111101100010100000000;
filter5[8][382] = 35'b11111010111011001010101110001000000;
filter5[8][383] = 35'b11110111001001111001001000100000000;
filter5[8][384] = 35'b00000001000100111111111101010100000;
filter5[8][385] = 35'b11111111110001111011010110011100000;
filter5[8][386] = 35'b00000010110000001010001011000000000;
filter5[8][387] = 35'b00000001011010111011011001000110000;
filter5[8][388] = 35'b00000000100111101011000110111110000;
filter5[8][389] = 35'b00000100001111100011011100111000000;
filter5[8][390] = 35'b00000001001010001011110111111010000;
filter5[8][391] = 35'b11111111100000010011101010111100100;
filter5[8][392] = 35'b11111011010100100010000111000000000;
filter5[8][393] = 35'b11111110101000110111101110111110000;
filter5[8][394] = 35'b11111111101100110010000100101001000;
filter5[8][395] = 35'b00000010101101000010111101011000000;
filter5[8][396] = 35'b00000010000111111011110011110100000;
filter5[8][397] = 35'b00000001101001111001110100111100000;
filter5[8][398] = 35'b00000010000010001010001111101000000;
filter5[8][399] = 35'b00000011000001101100000000001100000;
filter5[8][400] = 35'b00000010011101001000100001001100000;
filter5[8][401] = 35'b00000001011111111111011011110010000;
filter5[8][402] = 35'b11111111011100010101100111100110000;
filter5[8][403] = 35'b00000000001011001010110111011101000;
filter5[8][404] = 35'b00000011011100101000010011000000000;
filter5[8][405] = 35'b00000000000011111110111101001000011;
filter5[8][406] = 35'b11111101111001111010001000100100000;
filter5[8][407] = 35'b00000000000100101001001011100010101;
filter5[8][408] = 35'b00000000100111000110101001000111000;
filter5[8][409] = 35'b00000010110110011011100111000000000;
filter5[8][410] = 35'b00000001110101011111100101001000000;
filter5[8][411] = 35'b11111111110001000011111011011000010;
filter5[8][412] = 35'b00000001110100011100111011000100000;
filter5[8][413] = 35'b00000000111100110001001001111101000;
filter5[8][414] = 35'b00000001000001001001111110101000000;
filter5[8][415] = 35'b11111101111111111101011100100000000;
filter5[8][416] = 35'b11111110111000100000101100000100000;
filter5[8][417] = 35'b00000000000001111100011101000001111;
filter5[8][418] = 35'b11111110111110011100010101010000000;
filter5[8][419] = 35'b00000010001110000111100000100000000;
filter5[8][420] = 35'b00000000010100101111110100100101000;
filter5[8][421] = 35'b11111111110110101010011000011001000;
filter5[8][422] = 35'b11111111001110000110000111101001000;
filter5[8][423] = 35'b11111101101111001011100011001100000;
filter5[8][424] = 35'b00000010011000100010010011100100000;
filter5[8][425] = 35'b11111111111111100011010010100010111;
filter5[8][426] = 35'b11111100100011000011011011111100000;
filter5[8][427] = 35'b11111100101001111010001000010000000;
filter5[8][428] = 35'b11111100110001100101100010111000000;
filter5[8][429] = 35'b00000011100100110000001110110100000;
filter5[8][430] = 35'b11111100111101000000011100011000000;
filter5[8][431] = 35'b00000000101001010111101111000001000;
filter5[8][432] = 35'b11111110011111111111011110100000000;
filter5[8][433] = 35'b11111111000110100010110000011010000;
filter5[8][434] = 35'b11111111100010011000101100111111100;
filter5[8][435] = 35'b11011110111100001100111110000000000;
filter5[8][436] = 35'b11111000001011010100001011100000000;
filter5[8][437] = 35'b11110111111001011010100000110000000;
filter5[8][438] = 35'b00000000011111111101101111011111000;
filter5[8][439] = 35'b00000010001000111011000001011100000;
filter5[8][440] = 35'b11111111011011111010111100111011000;
filter5[8][441] = 35'b00000111110011100110010111100000000;
filter5[8][442] = 35'b00000001001011100111001000010010000;
filter5[8][443] = 35'b11111011101100111101010011010000000;
filter5[8][444] = 35'b11111111010100000001110011001010000;
filter5[8][445] = 35'b11111110101010111111111001111100000;
filter5[8][446] = 35'b00000001010000000010101000010000000;
filter5[8][447] = 35'b00000010110110000101011110000000000;
filter5[8][448] = 35'b11111111110110010110001100100100100;
filter5[8][449] = 35'b00000100110100001110100011101000000;
filter5[8][450] = 35'b11111011110000101100001101000000000;
filter5[8][451] = 35'b11111110110010001101101100111010000;
filter5[8][452] = 35'b11111010100111010101001101010000000;
filter5[8][453] = 35'b00000101101101100101001101110000000;
filter5[8][454] = 35'b11111101010110101011010000010100000;
filter5[8][455] = 35'b11111100101110101110100010100000000;
filter5[8][456] = 35'b00000000010101001011010110001000000;
filter5[8][457] = 35'b00000001000100010000110101011110000;
filter5[8][458] = 35'b00000011001100100000010010000000000;
filter5[8][459] = 35'b11111100000100001101101111000100000;
filter5[8][460] = 35'b00000000101101101001101001100100000;
filter5[8][461] = 35'b11111011101100011101010100101000000;
filter5[8][462] = 35'b00000001100101111001100000010110000;
filter5[8][463] = 35'b00000001000101011010110011110100000;
filter5[8][464] = 35'b00000100000001100011101010001000000;
filter5[8][465] = 35'b00000000101110111001101011001111000;
filter5[8][466] = 35'b11111111100000101110000001111101100;
filter5[8][467] = 35'b11111101010111101111111000000000000;
filter5[8][468] = 35'b00000101111011000110001011000000000;
filter5[8][469] = 35'b00000011010011010111011011110100000;
filter5[8][470] = 35'b11111001101100111000000011010000000;
filter5[8][471] = 35'b11111110111000000010101101111010000;
filter5[8][472] = 35'b00000010110110111000010111110000000;
filter5[8][473] = 35'b00000011110101110001110011111100000;
filter5[8][474] = 35'b11111110111001111111001110110100000;
filter5[8][475] = 35'b11110111100101010101010000100000000;
filter5[8][476] = 35'b00000000011101011011100001110000100;
filter5[8][477] = 35'b11111100000110001011110111100000000;
filter5[8][478] = 35'b11111101101001101010001101010100000;
filter5[8][479] = 35'b11111111110101110100101110110000110;
filter5[8][480] = 35'b11111001100011001110000001010000000;
filter5[8][481] = 35'b11111111100011110001011100100011000;
filter5[8][482] = 35'b11111101110001100100000001110000000;
filter5[8][483] = 35'b11111111000100100110101010100110000;
filter5[8][484] = 35'b11111001101001111100001111101000000;
filter5[8][485] = 35'b11111011011110101001011111011000000;
filter5[8][486] = 35'b11111001100100010001110100001000000;
filter5[8][487] = 35'b11111011001001011111011101011000000;
filter5[8][488] = 35'b11111101001100001100011111000000000;
filter5[8][489] = 35'b11111011101111101011111001011000000;
filter5[8][490] = 35'b11111000001001011110001000010000000;
filter5[8][491] = 35'b11111111010011111000011110010101000;
filter5[8][492] = 35'b11111010000010010001100000101000000;
filter5[8][493] = 35'b11110110010110000111011110000000000;
filter5[8][494] = 35'b11111100100100110001010110110100000;
filter5[8][495] = 35'b11111110100000001110000110010100000;
filter5[8][496] = 35'b11111100100111100010110000001100000;
filter5[8][497] = 35'b00000000011001100110100101000011100;
filter5[8][498] = 35'b11111100011100011111110110111100000;
filter5[8][499] = 35'b11111111111100111000101001000100101;
filter5[8][500] = 35'b00000101001011110000101101010000000;
filter5[8][501] = 35'b00000001000001000001110000100110000;
filter5[8][502] = 35'b11111110111011001011010001010110000;
filter5[8][503] = 35'b11111101110000001111001101000000000;
filter5[8][504] = 35'b11111111010100011011110111110010000;
filter5[8][505] = 35'b00000011100000110101100100111000000;
filter5[8][506] = 35'b00000001101010101110000100111000000;
filter5[8][507] = 35'b11111111111001111100010001000101110;
filter5[8][508] = 35'b11111011010101010011000000011000000;
filter5[8][509] = 35'b00000111001000101111010111100000000;
filter5[8][510] = 35'b00000011010001110010010001101000000;
filter5[8][511] = 35'b00000000100110010001101111110100000;
filter5[8][512] = 35'b11111110101100101010000111011100000;
filter5[8][513] = 35'b11111100100001100111100001110100000;
filter5[8][514] = 35'b00000000111010001001001110100000000;
filter5[8][515] = 35'b00000001011100000111110110001010000;
filter5[8][516] = 35'b00000001100011011000010010001000000;
filter5[8][517] = 35'b00000011110000100110001101100000000;
filter5[8][518] = 35'b11111101001111110000001001011100000;
filter5[8][519] = 35'b00000010110011010111010001100000000;
filter5[8][520] = 35'b11111101000110111000011100011100000;
filter5[8][521] = 35'b00000010000110010001001100110000000;
filter5[8][522] = 35'b11111110000111000000111101000010000;
filter5[8][523] = 35'b00000110001010110011010001010000000;
filter5[8][524] = 35'b11111110110011010111011110000010000;
filter5[8][525] = 35'b00000001000111110110010001001010000;
filter5[8][526] = 35'b00000111100101010101101000100000000;
filter5[8][527] = 35'b00000001100110001000001000001110000;
filter5[8][528] = 35'b11111110111111001010001011001100000;
filter5[8][529] = 35'b00000010011111011110111011111000000;
filter5[8][530] = 35'b00000011110000010100111001110100000;
filter5[8][531] = 35'b00000000011111111100000001100011000;
filter5[8][532] = 35'b00000000111000011010010100010100000;
filter5[8][533] = 35'b00000100110000010011100101010000000;
filter5[8][534] = 35'b00000001000110110001111010011000000;
filter5[8][535] = 35'b11111101101110011001000110011100000;
filter5[8][536] = 35'b11111111111101101110111110111100100;
filter5[8][537] = 35'b00000000010000110100110101100101000;
filter5[8][538] = 35'b11111111100110010010111010001000100;
filter5[8][539] = 35'b00000001101101110101100001110000000;
filter5[8][540] = 35'b00000001000001100000010111100010000;
filter5[8][541] = 35'b00000000011101101001100101000101000;
filter5[8][542] = 35'b11111110110111101101011011000110000;
filter5[8][543] = 35'b11111111000010010011011101010110000;
filter5[8][544] = 35'b11111111000010110000111000100111000;
filter5[8][545] = 35'b00000000100011101101000101100111000;
filter5[8][546] = 35'b11111110011001000111001010110000000;
filter5[8][547] = 35'b00000000000110001011010001111111000;
filter5[8][548] = 35'b11111100110001001101011111100100000;
filter5[8][549] = 35'b00000000011001011011111100011110100;
filter5[8][550] = 35'b11111110000111111100001110011110000;
filter5[8][551] = 35'b11111111000100000100011110111100000;
filter5[8][552] = 35'b00000001111110110001000011001100000;
filter5[8][553] = 35'b00000001010111011010010010011000000;
filter5[8][554] = 35'b00000001100010110000111001001110000;
filter5[8][555] = 35'b00000100010100010111000001101000000;
filter5[8][556] = 35'b11111011010000000000111000111000000;
filter5[8][557] = 35'b00000000101110100100000111111111000;
filter5[8][558] = 35'b00000010110011101101010010001000000;
filter5[8][559] = 35'b11111111000110110100110011000100000;
filter5[8][560] = 35'b11111111101101000100011000100000100;
filter5[8][561] = 35'b11111111011011001110110000000101000;
filter5[8][562] = 35'b11111110011111110100110100100010000;
filter5[8][563] = 35'b00000010111111101110111101010000000;
filter5[8][564] = 35'b11111100010011011010000010001100000;
filter5[8][565] = 35'b00000001000011110011011010000000000;
filter5[8][566] = 35'b11111100101000000000010111001000000;
filter5[8][567] = 35'b00000010000100111001110010011000000;
filter5[8][568] = 35'b11111110101010001000111001000010000;
filter5[8][569] = 35'b11111101000001010100010011110100000;
filter5[8][570] = 35'b11111101001101110101101000110100000;
filter5[8][571] = 35'b00000011000011000010111101010000000;
filter5[8][572] = 35'b11111101100001101001110110101100000;
filter5[8][573] = 35'b00000001001101101111010101110000000;
filter5[8][574] = 35'b11111100010111101011010111000000000;
filter5[8][575] = 35'b00000101000110001010011000101000000;
filter5[8][576] = 35'b00000000111001011011000101001101000;
filter5[8][577] = 35'b11111101100010001000011110001000000;
filter5[8][578] = 35'b00000000001011010111001000010110000;
filter5[8][579] = 35'b00000100101011010100010110101000000;
filter5[8][580] = 35'b00000011110111111100010100101000000;
filter5[8][581] = 35'b00000010100000010111100010110000000;
filter5[8][582] = 35'b11111111100010101011010011111101000;
filter5[8][583] = 35'b00000000000010110000010100011101011;
filter5[8][584] = 35'b11111101001000001010111010001000000;
filter5[8][585] = 35'b00000100100111111101110100101000000;
filter5[8][586] = 35'b00000000001111110010000101101000110;
filter5[8][587] = 35'b00000011111010000001110000110100000;
filter5[8][588] = 35'b00000010010111100101110000010000000;
filter5[8][589] = 35'b00000011001011100000100001110100000;
filter5[8][590] = 35'b00000001010101000100100000011100000;
filter5[8][591] = 35'b00000001110011010010101011101110000;
filter5[8][592] = 35'b00000001100000101101001001010010000;
filter5[8][593] = 35'b00000010001001101001100101001100000;
filter5[8][594] = 35'b00000001101100101011101100110000000;
filter5[8][595] = 35'b00000000111101010100001011000000000;
filter5[8][596] = 35'b11111111111110011111010010101011111;
filter5[8][597] = 35'b00000001100100011000110010000100000;
filter5[8][598] = 35'b11111110101110010101101110100100000;
filter5[8][599] = 35'b11111110010110110011100110010100000;
filter5[8][600] = 35'b11111100110111011000101111001100000;
filter5[8][601] = 35'b00000011111001100111101101101100000;
filter5[8][602] = 35'b11111101111001101000001101001000000;
filter5[8][603] = 35'b11111111111000111101010010111000101;
filter5[8][604] = 35'b11111110000000110110111011011110000;
filter5[8][605] = 35'b00000110001011011100110100011000000;
filter5[8][606] = 35'b11111110000011110001101001100100000;
filter5[8][607] = 35'b11111011010010111000000001100000000;
filter5[8][608] = 35'b11111111011001011101011010100011000;
filter5[8][609] = 35'b11111111101010110000110011110100000;
filter5[8][610] = 35'b11111001110110010010101010101000000;
filter5[8][611] = 35'b11111010001010111011100000100000000;
filter5[8][612] = 35'b00000011000100111001100101110000000;
filter5[8][613] = 35'b00000001000011010000010101101100000;
filter5[8][614] = 35'b11111110011000100001011011110000000;
filter5[8][615] = 35'b11111111111101110011110010100011000;
filter5[8][616] = 35'b11111111001000110101011100101000000;
filter5[8][617] = 35'b00000001000001010100100110001100000;
filter5[8][618] = 35'b00000011000100011010100100001100000;
filter5[8][619] = 35'b11111011010001000111001111001000000;
filter5[8][620] = 35'b11111011101100111000001111110000000;
filter5[8][621] = 35'b11111111110110110100000010111010110;
filter5[8][622] = 35'b00000001100111001000001010110100000;
filter5[8][623] = 35'b00000001111100001101010111011010000;
filter5[8][624] = 35'b00000001010011001001011000100110000;
filter5[8][625] = 35'b11111011010010101011010001011000000;
filter5[8][626] = 35'b00000000010100010001100101011010000;
filter5[8][627] = 35'b00000000101000110100111010000011000;
filter5[8][628] = 35'b11111101100110010011100100010100000;
filter5[8][629] = 35'b00000101111110101010001001111000000;
filter5[8][630] = 35'b11111100010001001111000100111000000;
filter5[8][631] = 35'b11111101010011111100101101100100000;
filter5[8][632] = 35'b00000010011000000100010011101000000;
filter5[8][633] = 35'b00000011000001001100001011010100000;
filter5[8][634] = 35'b11111111001111000111111010110101000;
filter5[8][635] = 35'b11111110011101110011010111100100000;
filter5[8][636] = 35'b00000010000001001101000000111000000;
filter5[8][637] = 35'b00000100100001011100101011010000000;
filter5[8][638] = 35'b11111001010101001001000101010000000;
filter5[8][639] = 35'b11111101111101101110001110101100000;
filter5[8][640] = 35'b11111110010110000101011011111100000;
filter5[8][641] = 35'b00000100000101111110001100011000000;
filter5[8][642] = 35'b11111110101010010110101100100010000;
filter5[8][643] = 35'b11111110000101000000011110000000000;
filter5[8][644] = 35'b11111010110110001101100100101000000;
filter5[8][645] = 35'b00000001101111111011110001110000000;
filter5[8][646] = 35'b11111110010111010011011000000010000;
filter5[8][647] = 35'b00000000001010001010011101110110110;
filter5[8][648] = 35'b00000000110110010101001100000101000;
filter5[8][649] = 35'b00000001000011101110001000011000000;
filter5[8][650] = 35'b11111111000110101110010110010001000;
filter5[8][651] = 35'b00000001100101100000110011101110000;
filter5[8][652] = 35'b00000010000110000011111010010000000;
filter5[8][653] = 35'b00000000000101011110101101100110011;
filter5[8][654] = 35'b00000100010100110101010001111000000;
filter5[8][655] = 35'b00000001111011110011000010110100000;
filter5[8][656] = 35'b11111101001010001100101101110100000;
filter5[8][657] = 35'b00000001000000100000101110011110000;
filter5[8][658] = 35'b11111011001110100110010010000000000;
filter5[8][659] = 35'b11110110110011011011010010000000000;
filter5[8][660] = 35'b00000100000011011000000001111000000;
filter5[8][661] = 35'b00000100010100010011010010000000000;
filter5[8][662] = 35'b00000011001101101010101110010100000;
filter5[8][663] = 35'b00000011010000000010100100110100000;
filter5[8][664] = 35'b00000010101011011000000101111100000;
filter5[8][665] = 35'b00000010100011001110110010110000000;
filter5[8][666] = 35'b11111010110000110011101011011000000;
filter5[8][667] = 35'b00000101010000101000101011110000000;
filter5[8][668] = 35'b11111111011010010001111100000101000;
filter5[8][669] = 35'b11111111010000110000110000011111000;
filter5[8][670] = 35'b11111111100000010110001000011100000;
filter5[8][671] = 35'b00000101000011001010000111001000000;
filter5[8][672] = 35'b11111111110101011010010010110000100;
filter5[8][673] = 35'b00000000011000100101001001101110100;
filter5[8][674] = 35'b00000000010000001101101000101100100;
filter5[8][675] = 35'b00000100011001000011101101101000000;
filter5[8][676] = 35'b00000000010001110101111111000100000;
filter5[8][677] = 35'b00000010110010011110111011001000000;
filter5[8][678] = 35'b11111101001010101000111001011000000;
filter5[8][679] = 35'b11111011001100010111110001010000000;
filter5[8][680] = 35'b00000001110010000101000111011010000;
filter5[8][681] = 35'b11111110100110010100101111100010000;
filter5[8][682] = 35'b11110110001101000110111110010000000;
filter5[8][683] = 35'b11111111001001010001000100000110000;
filter5[8][684] = 35'b11111000100000000000111001000000000;
filter5[8][685] = 35'b00000000101001011111100111000101000;
filter5[8][686] = 35'b00000000110000110000110010110000000;
filter5[8][687] = 35'b11111101110111001010101001101000000;
filter5[8][688] = 35'b00000001100011111001101011011110000;
filter5[8][689] = 35'b11111101101000111101100101110000000;
filter5[8][690] = 35'b11111011100001010101011001011000000;
filter5[8][691] = 35'b11111100010111010101110111011000000;
filter5[8][692] = 35'b11110111100101110100001010010000000;
filter5[8][693] = 35'b00000011001100110100001110100000000;
filter5[8][694] = 35'b11111111100110000110110001110010100;
filter5[8][695] = 35'b00000010001100100101111110100000000;
filter5[8][696] = 35'b00000011110000110111100011001100000;
filter5[8][697] = 35'b00000000001010000001110100010011110;
filter5[8][698] = 35'b00000011010110111010101001011000000;
filter5[8][699] = 35'b11111110000100000101110011001100000;
filter5[8][700] = 35'b11111101001110100110000010011100000;
filter5[8][701] = 35'b00000001100010000011100001010110000;
filter5[8][702] = 35'b00000001001110001000110001111100000;
filter5[8][703] = 35'b00000001000011110110111110011010000;
filter5[8][704] = 35'b11111111000100100010001101010010000;
filter5[8][705] = 35'b11111110111000111010011111101010000;
filter5[8][706] = 35'b11111110101011000001000111010110000;
filter5[8][707] = 35'b11111110111111010110000001011010000;
filter5[8][708] = 35'b11111110111000110110010011110010000;
filter5[8][709] = 35'b00000000001001111011111111100010110;
filter5[8][710] = 35'b00000000111011111000110101010110000;
filter5[8][711] = 35'b00000000111001000100011001101000000;
filter5[8][712] = 35'b11111111110000100010000010011001100;
filter5[8][713] = 35'b00000000011111101011000111111101000;
filter5[8][714] = 35'b11111111101001011000011111110011000;
filter5[8][715] = 35'b11111111010011100000000100101101000;
filter5[8][716] = 35'b11111110111110010010001101010100000;
filter5[8][717] = 35'b00000000010000110111011001100001100;
filter5[8][718] = 35'b11111111111000101011010111100100101;
filter5[8][719] = 35'b00000001000011011000111011110010000;
filter5[8][720] = 35'b00000000000001000000110111010001010;
filter5[8][721] = 35'b11111111101000011101111110001110100;
filter5[8][722] = 35'b00000000011101000010111001011000100;
filter5[8][723] = 35'b11111110000100100100100100100000000;
filter5[8][724] = 35'b00000000100011101011111000101001000;
filter5[8][725] = 35'b11111100100001100100010101000100000;
filter5[8][726] = 35'b00000000101001010110101110000001000;
filter5[8][727] = 35'b11111110111100011010111000001100000;
filter5[8][728] = 35'b11111110111000000010101010110010000;
filter5[8][729] = 35'b11111101111101100100011011101000000;
filter5[8][730] = 35'b11111010011101001110111111111000000;
filter5[8][731] = 35'b00000000101111010100011001010111000;
filter5[8][732] = 35'b11111110101010011100011010000010000;
filter5[8][733] = 35'b11111101110000011001001000111000000;
filter5[8][734] = 35'b00000000110111010110001011101000000;
filter5[8][735] = 35'b11111111001010101100011010101111000;
filter5[8][736] = 35'b11111110111100101000001101100010000;
filter5[8][737] = 35'b11111111000111010011000101010111000;
filter5[8][738] = 35'b11111011101100001010101000110000000;
filter5[8][739] = 35'b00000011000011110100111100111000000;
filter5[8][740] = 35'b11111011001001000010110111010000000;
filter5[8][741] = 35'b11111101001011011111100010000100000;
filter5[8][742] = 35'b11111100100001111001110010101100000;
filter5[8][743] = 35'b11111111010011101111101001111010000;
filter5[8][744] = 35'b11111011101111000010000111110000000;
filter5[8][745] = 35'b00000001000011001010000111101010000;
filter5[8][746] = 35'b00000001101100011100110111101000000;
filter5[8][747] = 35'b00000010101111011110010010100100000;
filter5[8][748] = 35'b11111111011100111000011010000110000;
filter5[8][749] = 35'b00000001010111100010001001010100000;
filter5[8][750] = 35'b11111010111111001010000101111000000;
filter5[8][751] = 35'b00000001010011111101000000101100000;
filter5[8][752] = 35'b11111100110110000001110001010000000;
filter5[8][753] = 35'b11111011001001001001110011000000000;
filter5[8][754] = 35'b00000011100001010111001110111100000;
filter5[8][755] = 35'b11111111001010111000110101101010000;
filter5[8][756] = 35'b11111111100101000000000001100011000;
filter5[8][757] = 35'b00000001100000001101011010000010000;
filter5[8][758] = 35'b00000001000011100101101101001100000;
filter5[8][759] = 35'b11111100000001101001100000110000000;
filter5[8][760] = 35'b11111111111110011101001100000111101;
filter5[8][761] = 35'b00000000011011001001100011100000100;
filter5[8][762] = 35'b00000010011100000000100000110000000;
filter5[8][763] = 35'b11111110100101001000100011010100000;
filter5[8][764] = 35'b00000000101111001101011111011110000;
filter5[8][765] = 35'b00000101000010110100110001100000000;
filter5[8][766] = 35'b00000000010001001110011100010010000;
filter5[8][767] = 35'b11111101110101101100110100111000000;
filter5[8][768] = 35'b11111111111000000000011010010110101;
filter5[8][769] = 35'b00000010010111100010010011101000000;
filter5[8][770] = 35'b11111111100010101000110000010000100;
filter5[8][771] = 35'b00000001111010111110010110010100000;
filter5[8][772] = 35'b11111111100101001011011010010110100;
filter5[8][773] = 35'b00000011011010010101010111011000000;
filter5[8][774] = 35'b11111101100101111001001011100000000;
filter5[8][775] = 35'b00000010110101010010010110110100000;
filter5[8][776] = 35'b00000001000100101100000101010000000;
filter5[8][777] = 35'b00000001101110000111000101010110000;
filter5[8][778] = 35'b00000011000010000000100111010100000;
filter5[8][779] = 35'b11111101111101110011010110000000000;
filter5[8][780] = 35'b00000001010101011101100101011010000;
filter5[8][781] = 35'b00000010100110000001110011001100000;
filter5[8][782] = 35'b00000101101011001000111010101000000;
filter5[8][783] = 35'b00000001100101010100111001001100000;
filter5[8][784] = 35'b00000011110111110111110110011100000;
filter5[8][785] = 35'b11111111100011000001001111010001000;
filter5[8][786] = 35'b11111101011111101001010011001000000;
filter5[8][787] = 35'b00000100101100100010100010100000000;
filter5[8][788] = 35'b11111010101110000101000011011000000;
filter5[8][789] = 35'b11111111000010010010100010111001000;
filter5[8][790] = 35'b00000001100111101011110011110000000;
filter5[8][791] = 35'b00000010001111100001111000011100000;
filter5[8][792] = 35'b11111111111000101000000000111000111;
filter5[8][793] = 35'b11111111011100111000101001101100000;
filter5[8][794] = 35'b00000011110111111011101000100100000;
filter5[8][795] = 35'b00000000100011100101110010111110000;
filter5[8][796] = 35'b11111111001010111111100100000001000;
filter5[8][797] = 35'b11111011101100100011011111001000000;
filter5[8][798] = 35'b11111100000110110101010000100000000;
filter5[8][799] = 35'b00000000000111001110010100000000100;
filter5[8][800] = 35'b00000000001110010101110111001001110;
filter5[8][801] = 35'b00000000001111101110100011011110110;
filter5[8][802] = 35'b11111111100011101001010100111101000;
filter5[8][803] = 35'b11111011111000000111010001110000000;
filter5[8][804] = 35'b00000100101101011100101100011000000;
filter5[8][805] = 35'b11111111110110100111110010000000100;
filter5[8][806] = 35'b11111110001101100011100110001100000;
filter5[8][807] = 35'b11111101010110101010010110000100000;
filter5[8][808] = 35'b11111111011111001010001000100101000;
filter5[8][809] = 35'b11111100011100110010010011010000000;
filter5[8][810] = 35'b00000000010011111100101001100001100;
filter5[8][811] = 35'b00000000101001101101111100001111000;
filter5[8][812] = 35'b00000000000000100000000110011110110;
filter5[8][813] = 35'b11111101110011001001000000101000000;
filter5[8][814] = 35'b11111011100000100111111111100000000;
filter5[8][815] = 35'b11111110111100100011101101111110000;
filter5[8][816] = 35'b11111111111011001010001100000010011;
filter5[8][817] = 35'b00000001001101111101110001110110000;
filter5[8][818] = 35'b11110100011010010110011001110000000;
filter5[8][819] = 35'b11111100100000111110111000101100000;
filter5[8][820] = 35'b11111101110110101011111101000000000;
filter5[8][821] = 35'b11111010110101100010011101000000000;
filter5[8][822] = 35'b11111111111100011100001111111100000;
filter5[8][823] = 35'b00000000111000110111110011011100000;
filter5[8][824] = 35'b11111101001000000010001010000100000;
filter5[8][825] = 35'b00000000110001110001001001010001000;
filter5[8][826] = 35'b00000101001111111111011001101000000;
filter5[8][827] = 35'b00000011101011001101001111001100000;
filter5[8][828] = 35'b11111100011001010011000010111000000;
filter5[8][829] = 35'b00000010001010010110010101111000000;
filter5[8][830] = 35'b00000011101100100001100000001100000;
filter5[8][831] = 35'b11111111100111100100100011111001000;
filter5[8][832] = 35'b11111111100100110100110101000110000;
filter5[8][833] = 35'b11111111111100011111010010110010011;
filter5[8][834] = 35'b11111111010101000001110101000110000;
filter5[8][835] = 35'b11111111111101010100100110000000001;
filter5[8][836] = 35'b11111110101111111110111111001010000;
filter5[8][837] = 35'b11111111111000100111001100101000010;
filter5[8][838] = 35'b00000000011101100101011110001010000;
filter5[8][839] = 35'b00000000001111000011110111110001110;
filter5[8][840] = 35'b00000000101000001001010011110100000;
filter5[8][841] = 35'b11111111101000000110101011100101100;
filter5[8][842] = 35'b11111111000011101010111010011011000;
filter5[8][843] = 35'b00000000010000010001101000100011100;
filter5[8][844] = 35'b11111111110100111011100111010010100;
filter5[8][845] = 35'b11111110110011001111101010100010000;
filter5[8][846] = 35'b00000000000111110000010111110000001;
filter5[8][847] = 35'b11111111100000010000001111010010100;
filter5[8][848] = 35'b11111111110011110101001000111000100;
filter5[8][849] = 35'b00000000010110010001001010011001000;
filter5[8][850] = 35'b11111110001010110110011001111010000;
filter5[8][851] = 35'b11111010000110001101000010101000000;
filter5[8][852] = 35'b11111101101011010110101111010000000;
filter5[8][853] = 35'b11111111010100101111010010100100000;
filter5[8][854] = 35'b11111110110011010111001101010100000;
filter5[8][855] = 35'b11111111111100101100111111100101110;
filter5[8][856] = 35'b00000000000001101111000110001001001;
filter5[8][857] = 35'b11111101101111001111110101011100000;
filter5[8][858] = 35'b11111100110110001110010011001000000;
filter5[8][859] = 35'b00000001000111111001000101001000000;
filter5[8][860] = 35'b11111111111010010111010111111111111;
filter5[8][861] = 35'b11111100100001101011010111111000000;
filter5[8][862] = 35'b00000001100011111001110110101110000;
filter5[8][863] = 35'b00000000101111100000100101110011000;
filter5[8][864] = 35'b11111101101000101011101110011100000;
filter5[8][865] = 35'b11111110000111011000010000010000000;
filter5[8][866] = 35'b11111100111001011011000101001000000;
filter5[8][867] = 35'b11111100001100101100001100011100000;
filter5[8][868] = 35'b11111111001110000101010111010010000;
filter5[8][869] = 35'b00000000000101010000100000101111111;
filter5[8][870] = 35'b11111110110111010100010100000010000;
filter5[8][871] = 35'b11111111010011100001011101100110000;
filter5[8][872] = 35'b11111101011110011000010010010000000;
filter5[8][873] = 35'b00000010111000111011100101100100000;
filter5[8][874] = 35'b00000000001010101001000000101011110;
filter5[8][875] = 35'b11111101111011000110111000010000000;
filter5[8][876] = 35'b00000000011111011011110000010011000;
filter5[8][877] = 35'b11111101000011001010010001111000000;
filter5[8][878] = 35'b11111111000011011001111111100011000;
filter5[8][879] = 35'b11111101111100111100101001100000000;
filter5[8][880] = 35'b11111101010010100100111010101000000;
filter5[8][881] = 35'b11111100000110001000100000011000000;
filter5[8][882] = 35'b00000011000011110001110100111000000;
filter5[8][883] = 35'b11111110110110101000000111110010000;
filter5[8][884] = 35'b00000000010100100010110001101100100;
filter5[8][885] = 35'b00001000000001100111011011100000000;
filter5[8][886] = 35'b00000001011100111100010010010010000;
filter5[8][887] = 35'b11111101000101100001101111000000000;
filter5[8][888] = 35'b00000001010011110100100101110000000;
filter5[8][889] = 35'b11111111011011010110101110111000000;
filter5[8][890] = 35'b11111111000100010110000001110001000;
filter5[8][891] = 35'b00000000001011000110011001110110100;
filter5[8][892] = 35'b11111111100110100011100111011011100;
filter5[8][893] = 35'b00000100011001001011001000000000000;
filter5[8][894] = 35'b11111011101100101101100100010000000;
filter5[8][895] = 35'b00000000101000101010110101001001000;
filter5[8][896] = 35'b11111110101010001111001010100000000;
filter5[8][897] = 35'b00000001100110101001110001101010000;
filter5[8][898] = 35'b00000100110101111010110011011000000;
filter5[8][899] = 35'b00000000111101011101110001011010000;
filter5[8][900] = 35'b11110011100100100110001001010000000;
filter5[8][901] = 35'b11111111010110101111010011000011000;
filter5[8][902] = 35'b11111110000001100001000111111010000;
filter5[8][903] = 35'b00000110101000101100100010011000000;
filter5[8][904] = 35'b00000001000111100000000100000100000;
filter5[8][905] = 35'b11111101111010101100000001001000000;
filter5[8][906] = 35'b00000010011100000111001010100100000;
filter5[8][907] = 35'b11111101110001010011010010011100000;
filter5[8][908] = 35'b00000001011111010100001010110110000;
filter5[8][909] = 35'b11111100001001001100111111100100000;
filter5[8][910] = 35'b00000010011001101100010001010000000;
filter5[8][911] = 35'b11111010000001100000001011000000000;
filter5[8][912] = 35'b11111101110000000010110000011000000;
filter5[8][913] = 35'b11111111010001000100001001110010000;
filter5[8][914] = 35'b11110010001100001110110001000000000;
filter5[8][915] = 35'b00000110101000111100110111101000000;
filter5[8][916] = 35'b00000100101001001100111101001000000;
filter5[8][917] = 35'b11110000001111110010100101100000000;
filter5[8][918] = 35'b11110110001011000011011010010000000;
filter5[8][919] = 35'b11111011010100111000110000111000000;
filter5[8][920] = 35'b11111110101000101100101110010000000;
filter5[8][921] = 35'b11111001010001001111101000001000000;
filter5[8][922] = 35'b11111001111100001010101001000000000;
filter5[8][923] = 35'b00000000111010001101001100101011000;
filter5[8][924] = 35'b00000010001111011011110000001000000;
filter5[8][925] = 35'b11110110100101001101001000010000000;
filter5[8][926] = 35'b00000001010111001110110110110000000;
filter5[8][927] = 35'b11111010001101001101000011000000000;
filter5[8][928] = 35'b00000001000110100000110111101010000;
filter5[8][929] = 35'b11110111000011011001100000010000000;
filter5[8][930] = 35'b11111100101111010000000001110100000;
filter5[8][931] = 35'b11111011000010011110010100111000000;
filter5[8][932] = 35'b11111101010010101011011010010100000;
filter5[8][933] = 35'b11111111101110111111100010101101100;
filter5[8][934] = 35'b11111110000111110001100111011100000;
filter5[8][935] = 35'b11111010000000110001010110000000000;
filter5[8][936] = 35'b11111010011000110101011111001000000;
filter5[8][937] = 35'b00000010100011100011010000111000000;
filter5[8][938] = 35'b00000001110101001001000111101100000;
filter5[8][939] = 35'b00000001100010101000000100011100000;
filter5[8][940] = 35'b00000001011101011011111000101110000;
filter5[8][941] = 35'b11111100000110111010001101110100000;
filter5[8][942] = 35'b11111010110000000100011001010000000;
filter5[8][943] = 35'b11101111101111011000000100100000000;
filter5[8][944] = 35'b11111101101111001100010010111000000;
filter5[8][945] = 35'b11111100001100011010110001000100000;
filter5[8][946] = 35'b00000001111100010100011101101000000;
filter5[8][947] = 35'b11111111010111100110110101110101000;
filter5[8][948] = 35'b11111111100111101100010010010100100;
filter5[8][949] = 35'b00000011110100011000100111011000000;
filter5[8][950] = 35'b00001001101000101111011000100000000;
filter5[8][951] = 35'b11111101111000011101111010100000000;
filter5[8][952] = 35'b11111101011010010010001110011100000;
filter5[8][953] = 35'b11110101001010100001110001000000000;
filter5[8][954] = 35'b11111100001101000110101001111100000;
filter5[8][955] = 35'b00000001110000100111010001110000000;
filter5[8][956] = 35'b00000101011110110000001000011000000;
filter5[8][957] = 35'b00000111001110000111000001010000000;
filter5[8][958] = 35'b11100111101110000011010000100000000;
filter5[8][959] = 35'b11111011000110111010110101001000000;
filter5[8][960] = 35'b00000101111000010100111111101000000;
filter5[8][961] = 35'b00000110100001110001101101111000000;
filter5[8][962] = 35'b00000000000110100111100111010000001;
filter5[8][963] = 35'b00000101111001100101101100011000000;
filter5[8][964] = 35'b11111011000110111010000101000000000;
filter5[8][965] = 35'b00000010111000001001100010110000000;
filter5[8][966] = 35'b00000011100100001110110000101100000;
filter5[8][967] = 35'b00000001111010000101001100100100000;
filter5[8][968] = 35'b00000010111001010101111110101100000;
filter5[8][969] = 35'b00001001011111011001001101000000000;
filter5[8][970] = 35'b11111111110011011001000100000001100;
filter5[8][971] = 35'b11111011011011111101000110000000000;
filter5[8][972] = 35'b11111011001110100101100100101000000;
filter5[8][973] = 35'b11111010000010111110100011101000000;
filter5[8][974] = 35'b00000001101010110010111101000000000;
filter5[8][975] = 35'b00000110111011001111000101010000000;
filter5[8][976] = 35'b11111110100010110010010010101110000;
filter5[8][977] = 35'b00000000000111110011111011101000010;
filter5[8][978] = 35'b11111110010110101101100100001110000;
filter5[8][979] = 35'b11111010000010100000111101110000000;
filter5[8][980] = 35'b00000011110000111111100010100100000;
filter5[8][981] = 35'b11111111001011111010011011001010000;
filter5[8][982] = 35'b11110100001111110111011011000000000;
filter5[8][983] = 35'b11110101011000010010011000110000000;
filter5[8][984] = 35'b00000001010101101000110111000100000;
filter5[8][985] = 35'b11111100111010001110100000100000000;
filter5[8][986] = 35'b11110111010000000001011011000000000;
filter5[8][987] = 35'b11111110101011000010111011010000000;
filter5[8][988] = 35'b00000010000011010101100000110100000;
filter5[8][989] = 35'b00000011100101100110101000000100000;
filter5[8][990] = 35'b00000000101111011011110000110111000;
filter5[8][991] = 35'b00000011111100111000100111000100000;
filter5[8][992] = 35'b11111100100011001000000010110100000;
filter5[8][993] = 35'b00000000110000101100011111000101000;
filter5[8][994] = 35'b11111101011011110000001011000100000;
filter5[8][995] = 35'b00000000101010100010110111110000000;
filter5[8][996] = 35'b11111011101011010010000110110000000;
filter5[8][997] = 35'b00000010101101001001101100111100000;
filter5[8][998] = 35'b11111101110100011001101010010100000;
filter5[8][999] = 35'b11111100100101011000101100011100000;
filter5[8][1000] = 35'b11111011100101110001110111100000000;
filter5[8][1001] = 35'b11111000001111011011100000100000000;
filter5[8][1002] = 35'b11111111010000110000000000101110000;
filter5[8][1003] = 35'b00000100110100001001001101010000000;
filter5[8][1004] = 35'b11111100011111001100111100101100000;
filter5[8][1005] = 35'b00000100000100001111100001000000000;
filter5[8][1006] = 35'b00000010001111001010100100010000000;
filter5[8][1007] = 35'b11111111010110101011011011110000000;
filter5[8][1008] = 35'b00000000101100010100101000111011000;
filter5[8][1009] = 35'b00000100010000000011000011110000000;
filter5[8][1010] = 35'b11111011010001010001100011100000000;
filter5[8][1011] = 35'b00000011100010001110111000110000000;
filter5[8][1012] = 35'b11111001011100100111010000011000000;
filter5[8][1013] = 35'b00001101001101010010101110110000000;
filter5[8][1014] = 35'b11111001111011111000011000110000000;
filter5[8][1015] = 35'b11111010011110100000001000000000000;
filter5[8][1016] = 35'b11111011100110100010001110011000000;
filter5[8][1017] = 35'b00000000000111001101011000001110010;
filter5[8][1018] = 35'b11101011100110100011101100000000000;
filter5[8][1019] = 35'b11111111100000111110101011000101100;
filter5[8][1020] = 35'b00000110100111111100000111011000000;
filter5[8][1021] = 35'b11111111111011100111011011101110010;
filter5[8][1022] = 35'b11110000010010100011011001000000000;
filter5[8][1023] = 35'b11111100010001000000110000110100000;
filter5[9][0] = 35'b11111111100111100010110001000101100;
filter5[9][1] = 35'b11111011111001111110100100110000000;
filter5[9][2] = 35'b11111110110101010111100101000100000;
filter5[9][3] = 35'b00000101011011000011111011010000000;
filter5[9][4] = 35'b00000000101101000000101001000000000;
filter5[9][5] = 35'b11111010001001100010001100010000000;
filter5[9][6] = 35'b11111111010110001111100101111000000;
filter5[9][7] = 35'b11111011000111010010101010001000000;
filter5[9][8] = 35'b00000001101101000100100001011010000;
filter5[9][9] = 35'b00000110001000001010110011001000000;
filter5[9][10] = 35'b11111100000101001010011001111000000;
filter5[9][11] = 35'b00000011110101000110110101001100000;
filter5[9][12] = 35'b00000011101011000100100000000000000;
filter5[9][13] = 35'b11111011110010000110100101011000000;
filter5[9][14] = 35'b11111101001101100111101011100100000;
filter5[9][15] = 35'b00000000111010011001101101011100000;
filter5[9][16] = 35'b11111111110010001011011100111101110;
filter5[9][17] = 35'b11111101100111000011101000100100000;
filter5[9][18] = 35'b00000011011101100001111010011100000;
filter5[9][19] = 35'b11111101111011010011100011001000000;
filter5[9][20] = 35'b11111101001101001110101100110000000;
filter5[9][21] = 35'b11111110001101111101100000100110000;
filter5[9][22] = 35'b11111100111011000001110100100100000;
filter5[9][23] = 35'b11111010010110000110100011110000000;
filter5[9][24] = 35'b11111111010100101001110101110101000;
filter5[9][25] = 35'b11111111000000010001001110100100000;
filter5[9][26] = 35'b11111111110101001111100101100010010;
filter5[9][27] = 35'b00000001001100011011101111001100000;
filter5[9][28] = 35'b00000001101001001110000101001010000;
filter5[9][29] = 35'b11111100011111001101100000111000000;
filter5[9][30] = 35'b00000100110101011010011010011000000;
filter5[9][31] = 35'b11110101111100010110011010010000000;
filter5[9][32] = 35'b11111101011101011001100001000000000;
filter5[9][33] = 35'b11111010100010011001100101111000000;
filter5[9][34] = 35'b00000001011101011000010110010100000;
filter5[9][35] = 35'b11111110110100010110110011001110000;
filter5[9][36] = 35'b11111110111110010100110000101010000;
filter5[9][37] = 35'b11111110110101000001100110001010000;
filter5[9][38] = 35'b00000110111100000010111111001000000;
filter5[9][39] = 35'b00000101100000000000011101101000000;
filter5[9][40] = 35'b00000000100010111111111111101110000;
filter5[9][41] = 35'b11111111001010000001101001110001000;
filter5[9][42] = 35'b00000000100110010100110010101101000;
filter5[9][43] = 35'b11111110100110001101101100001110000;
filter5[9][44] = 35'b00000010101000010001111101010000000;
filter5[9][45] = 35'b00000001111011010111111111101010000;
filter5[9][46] = 35'b00001100100101101110111100110000000;
filter5[9][47] = 35'b11111001110110100011110000000000000;
filter5[9][48] = 35'b11111110010011001000001101011100000;
filter5[9][49] = 35'b00000001111100100000011110001100000;
filter5[9][50] = 35'b11111111001111010001111101110010000;
filter5[9][51] = 35'b11111110011101010011010011011010000;
filter5[9][52] = 35'b11111111100000100100100100100111100;
filter5[9][53] = 35'b00000010001100000101001100010100000;
filter5[9][54] = 35'b00000011010101100100111110010100000;
filter5[9][55] = 35'b00000000100101111000010011100110000;
filter5[9][56] = 35'b00000101111110101010110010100000000;
filter5[9][57] = 35'b11111101101001101110111110011000000;
filter5[9][58] = 35'b11111111000101011111010100000111000;
filter5[9][59] = 35'b11111111101101010010001000001111100;
filter5[9][60] = 35'b00000000010100011010111000111010100;
filter5[9][61] = 35'b11111001111111001000110111001000000;
filter5[9][62] = 35'b11111110001011111100000001100110000;
filter5[9][63] = 35'b00000100110001001001110110100000000;
filter5[9][64] = 35'b11111100101010011110100001011000000;
filter5[9][65] = 35'b00000001100001111100101111010100000;
filter5[9][66] = 35'b11111110011100111000011110011000000;
filter5[9][67] = 35'b11111110111110110100110011100000000;
filter5[9][68] = 35'b11111110011011101111001000010010000;
filter5[9][69] = 35'b00000001000110000100000001010010000;
filter5[9][70] = 35'b00000000100111100000100000000101000;
filter5[9][71] = 35'b00000000001001011011000010111100110;
filter5[9][72] = 35'b00000000011110111001000110111011100;
filter5[9][73] = 35'b00000010001010110011000100000100000;
filter5[9][74] = 35'b11111110011000101000011000001000000;
filter5[9][75] = 35'b00000001011100010110110000111000000;
filter5[9][76] = 35'b00000001111001100011010101010000000;
filter5[9][77] = 35'b11111111110001010110100100111111000;
filter5[9][78] = 35'b00000000110010111010001001001100000;
filter5[9][79] = 35'b11111101111111000110100011001000000;
filter5[9][80] = 35'b00000000101101001011010001011100000;
filter5[9][81] = 35'b00000000010101010101000001001000100;
filter5[9][82] = 35'b00000001011011111110101111011110000;
filter5[9][83] = 35'b11111111110101011110111101011000000;
filter5[9][84] = 35'b00000001111110101111011110100010000;
filter5[9][85] = 35'b11111111010100011110100000010100000;
filter5[9][86] = 35'b11111111110001101011001101110011010;
filter5[9][87] = 35'b11111111010101110000111001110101000;
filter5[9][88] = 35'b11111111101100010101001010101000000;
filter5[9][89] = 35'b00000000010100100010010101111001100;
filter5[9][90] = 35'b00000000101111011000111010000100000;
filter5[9][91] = 35'b11111111010011110110101000110000000;
filter5[9][92] = 35'b00000000111011101000001100101010000;
filter5[9][93] = 35'b11111110111001101111000101000110000;
filter5[9][94] = 35'b00000010000111011010100111111100000;
filter5[9][95] = 35'b11111101000010010101110101000000000;
filter5[9][96] = 35'b11111100101001011000000110111000000;
filter5[9][97] = 35'b11111110001010010011001011111010000;
filter5[9][98] = 35'b11111011100000100100000010100000000;
filter5[9][99] = 35'b11111100000110101100010101001000000;
filter5[9][100] = 35'b11111100011001110001111100000100000;
filter5[9][101] = 35'b00000001100000010110100110001010000;
filter5[9][102] = 35'b00000010111001010001011011001100000;
filter5[9][103] = 35'b00000100000101111000010010011000000;
filter5[9][104] = 35'b00000000110011101110101110000111000;
filter5[9][105] = 35'b00000011000000011011011111110000000;
filter5[9][106] = 35'b00000010001001110100011110010000000;
filter5[9][107] = 35'b11111110000111110111000100101010000;
filter5[9][108] = 35'b11111111011100001100010001101001000;
filter5[9][109] = 35'b11111110000001001100110100000010000;
filter5[9][110] = 35'b00000011100101101001111000110000000;
filter5[9][111] = 35'b00000111111101111001000101000000000;
filter5[9][112] = 35'b11111011100011101111011111111000000;
filter5[9][113] = 35'b00000000010101001001000110100000000;
filter5[9][114] = 35'b11111111001010010010111010010001000;
filter5[9][115] = 35'b00000111001001000100110101011000000;
filter5[9][116] = 35'b11111101100000011011111011011000000;
filter5[9][117] = 35'b11111001101010110101100101101000000;
filter5[9][118] = 35'b11111100111111001010110101110000000;
filter5[9][119] = 35'b00000001010011011100101010111100000;
filter5[9][120] = 35'b00000011011110011011101100101000000;
filter5[9][121] = 35'b11111111100111000101001000010100100;
filter5[9][122] = 35'b00000010011000111100010011101100000;
filter5[9][123] = 35'b00000100010101101010001100111000000;
filter5[9][124] = 35'b00000000101100011001110010100101000;
filter5[9][125] = 35'b11111001101100010100011010001000000;
filter5[9][126] = 35'b11111110001101011001111001111010000;
filter5[9][127] = 35'b11111110100000110011010100010100000;
filter5[9][128] = 35'b11110110011101111111101000000000000;
filter5[9][129] = 35'b11111000111100000111011111001000000;
filter5[9][130] = 35'b00000100100110111000101001000000000;
filter5[9][131] = 35'b11111001100000110001010000110000000;
filter5[9][132] = 35'b11110100010011101101010111100000000;
filter5[9][133] = 35'b11111011011000100101111010101000000;
filter5[9][134] = 35'b11111110000000100111110110010000000;
filter5[9][135] = 35'b11111111000101101101010111110010000;
filter5[9][136] = 35'b11111111101000100010111101100111100;
filter5[9][137] = 35'b11111111011100111000110011010100000;
filter5[9][138] = 35'b11101101101110110101010011100000000;
filter5[9][139] = 35'b11110100001011100110011001000000000;
filter5[9][140] = 35'b11111010100101001000011010011000000;
filter5[9][141] = 35'b11101000110000110111001011000000000;
filter5[9][142] = 35'b11110001100000110100101000010000000;
filter5[9][143] = 35'b11111101111011010100010010110100000;
filter5[9][144] = 35'b11111010111111000001011100000000000;
filter5[9][145] = 35'b11101000111110101101111100000000000;
filter5[9][146] = 35'b11110001011111100000111110100000000;
filter5[9][147] = 35'b11111111111100100101110001100011010;
filter5[9][148] = 35'b00000010011011111100101001010000000;
filter5[9][149] = 35'b11111101110011110001101101101000000;
filter5[9][150] = 35'b00000000100111110001111100101010000;
filter5[9][151] = 35'b00000010000111101101000111010000000;
filter5[9][152] = 35'b00000001101011110100001110101000000;
filter5[9][153] = 35'b00000110010011001010010010110000000;
filter5[9][154] = 35'b11111111011010111001000001011011000;
filter5[9][155] = 35'b11111111010011010001001000101101000;
filter5[9][156] = 35'b00000000001110001000000100110001010;
filter5[9][157] = 35'b11111111100010000111011011000110100;
filter5[9][158] = 35'b00000001000000010010101111111000000;
filter5[9][159] = 35'b00000001010110010111111100011110000;
filter5[9][160] = 35'b00000010010100011001111011010000000;
filter5[9][161] = 35'b11111010100010001110111011100000000;
filter5[9][162] = 35'b11111111010000010011011011101110000;
filter5[9][163] = 35'b11111100000000000000101001001100000;
filter5[9][164] = 35'b00000000100111111110100000010001000;
filter5[9][165] = 35'b11111111101110101001010101000001000;
filter5[9][166] = 35'b00000000111101011100011110000101000;
filter5[9][167] = 35'b00001000010010010010011101110000000;
filter5[9][168] = 35'b00001001111111000101011010100000000;
filter5[9][169] = 35'b00000010011000100010011011000000000;
filter5[9][170] = 35'b00000000010111001110111010010111000;
filter5[9][171] = 35'b11111110011101111111010010111000000;
filter5[9][172] = 35'b00000010110011001100010010000000000;
filter5[9][173] = 35'b11111101001001011001010100110000000;
filter5[9][174] = 35'b00000001010011011010010010001010000;
filter5[9][175] = 35'b00001100010000011011000001000000000;
filter5[9][176] = 35'b11110101010101111111110110100000000;
filter5[9][177] = 35'b11111011010010101111110010001000000;
filter5[9][178] = 35'b11111010010000111100110001000000000;
filter5[9][179] = 35'b00000010000000101001001101001000000;
filter5[9][180] = 35'b00000101111010000010111001110000000;
filter5[9][181] = 35'b11110110101000111111010111000000000;
filter5[9][182] = 35'b00001001110100000100111011000000000;
filter5[9][183] = 35'b00001001100110011001100101100000000;
filter5[9][184] = 35'b11110000000011001101010010100000000;
filter5[9][185] = 35'b11110010010101111010111000100000000;
filter5[9][186] = 35'b11101001111101001011011110000000000;
filter5[9][187] = 35'b11111100010000011001100110010100000;
filter5[9][188] = 35'b11110101001011100111110000110000000;
filter5[9][189] = 35'b11101101111011111100110101000000000;
filter5[9][190] = 35'b11111011011111101000101000100000000;
filter5[9][191] = 35'b11111011010001100101101110000000000;
filter5[9][192] = 35'b11111011101000100010101110000000000;
filter5[9][193] = 35'b11111010001101001111101110011000000;
filter5[9][194] = 35'b00000001110001110010101011100100000;
filter5[9][195] = 35'b11111011000101010010101011101000000;
filter5[9][196] = 35'b11111000110110010001001010111000000;
filter5[9][197] = 35'b00000010110110011010110010110100000;
filter5[9][198] = 35'b00000011110000101111000010011100000;
filter5[9][199] = 35'b00000010000101110110000110010100000;
filter5[9][200] = 35'b11110111011000010110001010000000000;
filter5[9][201] = 35'b11111110010011000000110010011110000;
filter5[9][202] = 35'b00000000011000110001000100000110100;
filter5[9][203] = 35'b11110110010101100000101011010000000;
filter5[9][204] = 35'b11111101000111100100100000110100000;
filter5[9][205] = 35'b11111101001100000100010001011100000;
filter5[9][206] = 35'b00000010111010011010010011011100000;
filter5[9][207] = 35'b11111110111110001110001110111100000;
filter5[9][208] = 35'b11111001101011110101101111101000000;
filter5[9][209] = 35'b11111011010001100010010001011000000;
filter5[9][210] = 35'b11110101000001110111010011110000000;
filter5[9][211] = 35'b11110001100110110011101010110000000;
filter5[9][212] = 35'b11111110101100100011100100001100000;
filter5[9][213] = 35'b11110100001010111101010101110000000;
filter5[9][214] = 35'b11111101111111101100000110111100000;
filter5[9][215] = 35'b11110000110111110101110010110000000;
filter5[9][216] = 35'b00010000000101001100010101100000000;
filter5[9][217] = 35'b00000110100001000100111100110000000;
filter5[9][218] = 35'b11110011101001111111010111000000000;
filter5[9][219] = 35'b11111111111111001110000100010100011;
filter5[9][220] = 35'b00000001000000000110111101110000000;
filter5[9][221] = 35'b00000011001100001001100101110000000;
filter5[9][222] = 35'b11111001011000010001111110111000000;
filter5[9][223] = 35'b11111110111110101010110100101000000;
filter5[9][224] = 35'b11101001100110011111100100100000000;
filter5[9][225] = 35'b11110111010110011010111010000000000;
filter5[9][226] = 35'b11111010001010010011001001111000000;
filter5[9][227] = 35'b11111100101111010000001100110100000;
filter5[9][228] = 35'b11111101010011010100111011011100000;
filter5[9][229] = 35'b00000001111101000001000110101000000;
filter5[9][230] = 35'b00000011111111000010001000101100000;
filter5[9][231] = 35'b00000000010010110100011101101101000;
filter5[9][232] = 35'b00001111000111100100011101000000000;
filter5[9][233] = 35'b11111100111111001000111000111100000;
filter5[9][234] = 35'b00000001010100010110110011011110000;
filter5[9][235] = 35'b00000011000101001100000110101100000;
filter5[9][236] = 35'b11111111001111010011010111000000000;
filter5[9][237] = 35'b11111011111001001001101011111000000;
filter5[9][238] = 35'b00000001111001001001111111110110000;
filter5[9][239] = 35'b00000001001011001101011110100010000;
filter5[9][240] = 35'b11111001000011111110110001101000000;
filter5[9][241] = 35'b11111111110011111001100001101100110;
filter5[9][242] = 35'b00000001111101011111001011000100000;
filter5[9][243] = 35'b11111101011000001100011101111100000;
filter5[9][244] = 35'b00000001100111011101110101110110000;
filter5[9][245] = 35'b11111110111100110011110011111110000;
filter5[9][246] = 35'b00000000001110111010100011011011110;
filter5[9][247] = 35'b00000000111010001101101000001101000;
filter5[9][248] = 35'b11110010001100000101010110110000000;
filter5[9][249] = 35'b11111101100100101010111110111100000;
filter5[9][250] = 35'b00000001111010001100011011110110000;
filter5[9][251] = 35'b00000100011100010110110101100000000;
filter5[9][252] = 35'b00000010111010000000001011100000000;
filter5[9][253] = 35'b11111001011010100101110100011000000;
filter5[9][254] = 35'b00000000100101101000100000101001000;
filter5[9][255] = 35'b11111100010100001101110101111100000;
filter5[9][256] = 35'b11111100111100011101100110101100000;
filter5[9][257] = 35'b00000000010111011100111010011011000;
filter5[9][258] = 35'b11111111000010001001011100101101000;
filter5[9][259] = 35'b11111100111010100011010101111100000;
filter5[9][260] = 35'b00000000000101000101110110010111010;
filter5[9][261] = 35'b11111110011111011110110100010100000;
filter5[9][262] = 35'b11111110111101110101111111100010000;
filter5[9][263] = 35'b00000010000110001110111011010100000;
filter5[9][264] = 35'b11111100111100001111110001000000000;
filter5[9][265] = 35'b11111111001111100011100000010000000;
filter5[9][266] = 35'b11111111111010001001111101001111011;
filter5[9][267] = 35'b00000001000100010110110110010100000;
filter5[9][268] = 35'b11111101010001000000101011111000000;
filter5[9][269] = 35'b11111110011010011000000011011010000;
filter5[9][270] = 35'b11111101100001101111011001000100000;
filter5[9][271] = 35'b11111100111110001101001001010000000;
filter5[9][272] = 35'b11111000010001011100101001100000000;
filter5[9][273] = 35'b11110110110100100110010000000000000;
filter5[9][274] = 35'b11101000001101111000011011100000000;
filter5[9][275] = 35'b11111001000000011000111110011000000;
filter5[9][276] = 35'b00000010101001110110100110011100000;
filter5[9][277] = 35'b11110101010001110011011101000000000;
filter5[9][278] = 35'b11101100101111110101110011100000000;
filter5[9][279] = 35'b11110101111110000100111001010000000;
filter5[9][280] = 35'b00001111010100000101000110000000000;
filter5[9][281] = 35'b11110110100111011110001010110000000;
filter5[9][282] = 35'b11111001111110100010101011100000000;
filter5[9][283] = 35'b00000011100100000010111110101100000;
filter5[9][284] = 35'b00001011011000011101100111110000000;
filter5[9][285] = 35'b11111000101110000100100010110000000;
filter5[9][286] = 35'b11111010000010000100000110111000000;
filter5[9][287] = 35'b11101110101101101010010000000000000;
filter5[9][288] = 35'b11110101110111100000000001110000000;
filter5[9][289] = 35'b11101001001001000000010010100000000;
filter5[9][290] = 35'b11111010010000010101001110100000000;
filter5[9][291] = 35'b11111100110000001010110011100100000;
filter5[9][292] = 35'b11111111000010100011000110111001000;
filter5[9][293] = 35'b11111010011001111111101001001000000;
filter5[9][294] = 35'b11111110110011001111000000011100000;
filter5[9][295] = 35'b00000011011011000100001001011000000;
filter5[9][296] = 35'b00001000001101010110000011000000000;
filter5[9][297] = 35'b00000010110101011110101101100100000;
filter5[9][298] = 35'b11111111001101010000000001000110000;
filter5[9][299] = 35'b00000011000101100000111101011000000;
filter5[9][300] = 35'b11111101010110111100010000100100000;
filter5[9][301] = 35'b11111111100010010100100011011100000;
filter5[9][302] = 35'b11111110010110101101100110010010000;
filter5[9][303] = 35'b11111110011101110100100001000100000;
filter5[9][304] = 35'b11101110000000000000010010100000000;
filter5[9][305] = 35'b00000001010000110011011001101000000;
filter5[9][306] = 35'b00000010110010010001111110101100000;
filter5[9][307] = 35'b11111111010110100000011111100101000;
filter5[9][308] = 35'b00000000010111000000100001101101000;
filter5[9][309] = 35'b11111110011001111100011110110010000;
filter5[9][310] = 35'b11111101111100000001100100011100000;
filter5[9][311] = 35'b11111001110100011001111000101000000;
filter5[9][312] = 35'b11110001000000001011110111100000000;
filter5[9][313] = 35'b11111111111010000010011010111010011;
filter5[9][314] = 35'b00000010111110001010101001111100000;
filter5[9][315] = 35'b00000000000010110110111011010101010;
filter5[9][316] = 35'b11111110110100000000111111000010000;
filter5[9][317] = 35'b11111011101110010001001010101000000;
filter5[9][318] = 35'b11110100111110101101011111010000000;
filter5[9][319] = 35'b00000011101000111010000000100000000;
filter5[9][320] = 35'b11111101110100110001111011110000000;
filter5[9][321] = 35'b11111100010101111101010111101000000;
filter5[9][322] = 35'b00000010010101101011100100000000000;
filter5[9][323] = 35'b11111010011100000101101010011000000;
filter5[9][324] = 35'b11111011101010100101111110110000000;
filter5[9][325] = 35'b00000000110000001001011010011011000;
filter5[9][326] = 35'b00000001111011101011001100110010000;
filter5[9][327] = 35'b00000111111101111010101000011000000;
filter5[9][328] = 35'b11111111110110001001101100011101010;
filter5[9][329] = 35'b11111110101101100010011011110010000;
filter5[9][330] = 35'b00000000001000010111010110100010110;
filter5[9][331] = 35'b11111110010011011011010111111000000;
filter5[9][332] = 35'b00000010000111101000101100110100000;
filter5[9][333] = 35'b11111010010010110000000010110000000;
filter5[9][334] = 35'b11111001010110111101010110000000000;
filter5[9][335] = 35'b00000010111111101110100010101100000;
filter5[9][336] = 35'b00000010110111111010111110010000000;
filter5[9][337] = 35'b11111100100111110000100000110000000;
filter5[9][338] = 35'b00000001000001010101000110001110000;
filter5[9][339] = 35'b11111110111101011111001010001110000;
filter5[9][340] = 35'b00000001001111101111000110010110000;
filter5[9][341] = 35'b11111110010010011111110011110000000;
filter5[9][342] = 35'b11111100001010001010111111011000000;
filter5[9][343] = 35'b11111101010000101011111010000100000;
filter5[9][344] = 35'b11111110111010001010111111010000000;
filter5[9][345] = 35'b11111110011011000100100111011110000;
filter5[9][346] = 35'b11111101001000000000001111001000000;
filter5[9][347] = 35'b11111110100100101001100001110100000;
filter5[9][348] = 35'b00000000011111011011110010010000000;
filter5[9][349] = 35'b11111110110011110101011100100000000;
filter5[9][350] = 35'b11111111010101100010011111101000000;
filter5[9][351] = 35'b11111100011101100110001011110100000;
filter5[9][352] = 35'b11111010110011011110101110000000000;
filter5[9][353] = 35'b11111011011100110100101000101000000;
filter5[9][354] = 35'b11111101010001010010001111010100000;
filter5[9][355] = 35'b00000001010101001010000110111110000;
filter5[9][356] = 35'b11111100010111100011110100111000000;
filter5[9][357] = 35'b11111100000101101111100101111100000;
filter5[9][358] = 35'b00000111010001100011110101110000000;
filter5[9][359] = 35'b00000101011100000101100101011000000;
filter5[9][360] = 35'b00000010110110101111010011110000000;
filter5[9][361] = 35'b11111111001001010101101000010000000;
filter5[9][362] = 35'b00000000111001101110100011010011000;
filter5[9][363] = 35'b11111110110001010101011111010000000;
filter5[9][364] = 35'b00000001011110101100000111111100000;
filter5[9][365] = 35'b11111100110010110111101111111100000;
filter5[9][366] = 35'b00000110110001010101111011100000000;
filter5[9][367] = 35'b11111011110001000110111100001000000;
filter5[9][368] = 35'b11111111001110100010000110010101000;
filter5[9][369] = 35'b11111110011001101110110111110100000;
filter5[9][370] = 35'b11111110110100010011101001101000000;
filter5[9][371] = 35'b00000011110000011011101101001100000;
filter5[9][372] = 35'b00000010111001101001100101110100000;
filter5[9][373] = 35'b11111100110101011101011110011100000;
filter5[9][374] = 35'b11111110110000101011100101001010000;
filter5[9][375] = 35'b00000010011010011110010010000000000;
filter5[9][376] = 35'b00000010001000110101110011010100000;
filter5[9][377] = 35'b00000001001010001010111000001000000;
filter5[9][378] = 35'b00000100000100111011110110001000000;
filter5[9][379] = 35'b11111110101111101110000110111110000;
filter5[9][380] = 35'b00000110001011011000101101000000000;
filter5[9][381] = 35'b11111010100110011110011111010000000;
filter5[9][382] = 35'b11111110011111101111101000111100000;
filter5[9][383] = 35'b11111110101100110100010010111010000;
filter5[9][384] = 35'b11111111100101100011101110110100100;
filter5[9][385] = 35'b00000010101100100101110000010100000;
filter5[9][386] = 35'b00000000000111111110011111010111100;
filter5[9][387] = 35'b11111110100101010001000001001100000;
filter5[9][388] = 35'b11111111101001000111010000010001100;
filter5[9][389] = 35'b00000000110001001011000111000111000;
filter5[9][390] = 35'b11111111001111010000111001101001000;
filter5[9][391] = 35'b11111110101011101110111111101110000;
filter5[9][392] = 35'b11111110101011100100101111110010000;
filter5[9][393] = 35'b00000010001001100111001101110100000;
filter5[9][394] = 35'b00000000010010101101010110011001000;
filter5[9][395] = 35'b11111111011001001110111010011011000;
filter5[9][396] = 35'b00000001100011011010011110010110000;
filter5[9][397] = 35'b11111111101100100001111100011100100;
filter5[9][398] = 35'b11111110010111100111001001100010000;
filter5[9][399] = 35'b00000011001100010001010000110000000;
filter5[9][400] = 35'b00000001001101100110011010000110000;
filter5[9][401] = 35'b11111110011110111010100110000010000;
filter5[9][402] = 35'b00000001000101100110100000101100000;
filter5[9][403] = 35'b00000000101001010111011111010011000;
filter5[9][404] = 35'b11111110101101011100001011000100000;
filter5[9][405] = 35'b11111101000011010111100010110000000;
filter5[9][406] = 35'b11111011101000101110101111010000000;
filter5[9][407] = 35'b00000000100100101011010000110101000;
filter5[9][408] = 35'b00000000111001111100111000110010000;
filter5[9][409] = 35'b00000000110111100010010110110100000;
filter5[9][410] = 35'b00000000011000111100111010101101000;
filter5[9][411] = 35'b11111110100011000110100011011000000;
filter5[9][412] = 35'b11111111001100011100100000001100000;
filter5[9][413] = 35'b11111111001110101101110101101000000;
filter5[9][414] = 35'b00000001100111001011110100111010000;
filter5[9][415] = 35'b00000001110000101011000000010000000;
filter5[9][416] = 35'b00000000100111101110110010011001000;
filter5[9][417] = 35'b11111111011110000011011010000110000;
filter5[9][418] = 35'b11111110111010010100101100011110000;
filter5[9][419] = 35'b11111110010101011100110101110100000;
filter5[9][420] = 35'b11111110111111010010110110001100000;
filter5[9][421] = 35'b00000000110011001110000110100111000;
filter5[9][422] = 35'b00000010010001011101111001111000000;
filter5[9][423] = 35'b00000010000111011001111111000100000;
filter5[9][424] = 35'b11111110011000000101101000000110000;
filter5[9][425] = 35'b11111111111010110111001010010111011;
filter5[9][426] = 35'b00000001110001001110011001110000000;
filter5[9][427] = 35'b11111111101001001000111110110110100;
filter5[9][428] = 35'b11111101110100011110000010010100000;
filter5[9][429] = 35'b11111101101011010001100101010000000;
filter5[9][430] = 35'b00000001101100010001110110000010000;
filter5[9][431] = 35'b11111111101000111100010100000011100;
filter5[9][432] = 35'b11111101110110001110001110001000000;
filter5[9][433] = 35'b00000001101110010110110100111110000;
filter5[9][434] = 35'b00000100011100011010101000111000000;
filter5[9][435] = 35'b11111000011101101010101111100000000;
filter5[9][436] = 35'b11111111110010011111010110011111110;
filter5[9][437] = 35'b11111111001011011101110101011110000;
filter5[9][438] = 35'b00000000101111100101010110111011000;
filter5[9][439] = 35'b11111100101001101111001101001100000;
filter5[9][440] = 35'b00000010100010100101000100100000000;
filter5[9][441] = 35'b00000010101010011111100011010000000;
filter5[9][442] = 35'b11111101110010010011000011001000000;
filter5[9][443] = 35'b11111000110101100110000110111000000;
filter5[9][444] = 35'b00000000100101011011101111011100000;
filter5[9][445] = 35'b00000010011010001001101011010000000;
filter5[9][446] = 35'b00000011001100000101100110000000000;
filter5[9][447] = 35'b00000101001110000001000111000000000;
filter5[9][448] = 35'b00000000010010110101100010011010100;
filter5[9][449] = 35'b11111100101001011111001001010100000;
filter5[9][450] = 35'b00000010001111000010001000001000000;
filter5[9][451] = 35'b11111101100011101100100111001100000;
filter5[9][452] = 35'b11111111101010001001010001111110000;
filter5[9][453] = 35'b00000011001001100110101100110100000;
filter5[9][454] = 35'b00000001101111010001110101110110000;
filter5[9][455] = 35'b11111101010010010000000010110000000;
filter5[9][456] = 35'b11111100100000000000000100101000000;
filter5[9][457] = 35'b00000100001011110101110001101000000;
filter5[9][458] = 35'b11111111011001100101011110011100000;
filter5[9][459] = 35'b11111101110000011010111101000100000;
filter5[9][460] = 35'b11111111011100011010100000000001000;
filter5[9][461] = 35'b00000010001000110001010110110100000;
filter5[9][462] = 35'b00000001100010010100000100111110000;
filter5[9][463] = 35'b00000101010000111010101011111000000;
filter5[9][464] = 35'b11111111000000100000010100000001000;
filter5[9][465] = 35'b11111111001011001100110101010010000;
filter5[9][466] = 35'b11111011011000110001011000001000000;
filter5[9][467] = 35'b11111111110010011001110100111101000;
filter5[9][468] = 35'b11111111110101110000100111001110010;
filter5[9][469] = 35'b00000000010111110101010010101010100;
filter5[9][470] = 35'b11111010111010011001111110001000000;
filter5[9][471] = 35'b11111111000101101111010000011000000;
filter5[9][472] = 35'b00000000111101111000010001111100000;
filter5[9][473] = 35'b00000110011110000110011100000000000;
filter5[9][474] = 35'b11111011111001011010011100011000000;
filter5[9][475] = 35'b11110111110010011101011010010000000;
filter5[9][476] = 35'b00000001100100000000110010010110000;
filter5[9][477] = 35'b00000100001101101010111001011000000;
filter5[9][478] = 35'b00000010100011101011010010010100000;
filter5[9][479] = 35'b11111100001001111110110000000000000;
filter5[9][480] = 35'b00000001111111100101111010001100000;
filter5[9][481] = 35'b00000010011000000000001111110000000;
filter5[9][482] = 35'b11111000101111101000100111100000000;
filter5[9][483] = 35'b11111111001001000111000011001111000;
filter5[9][484] = 35'b11111110000010000101100001101110000;
filter5[9][485] = 35'b11111010110111111001101000011000000;
filter5[9][486] = 35'b00000101010101000111010110010000000;
filter5[9][487] = 35'b00000001111000010010000011010100000;
filter5[9][488] = 35'b00000000011010111101111011100000100;
filter5[9][489] = 35'b00000000110110010000100101010000000;
filter5[9][490] = 35'b11101001100011100000000010100000000;
filter5[9][491] = 35'b11111101111111000011011001110000000;
filter5[9][492] = 35'b11111110000101101110010100011010000;
filter5[9][493] = 35'b11111110010010100100110111010100000;
filter5[9][494] = 35'b00000100010100001111011110000000000;
filter5[9][495] = 35'b00000111010000111110111101110000000;
filter5[9][496] = 35'b00000100011010000001011000011000000;
filter5[9][497] = 35'b11111111010011001101011101111101000;
filter5[9][498] = 35'b11111101101010100000011100010000000;
filter5[9][499] = 35'b11111011100010000100001101000000000;
filter5[9][500] = 35'b00000010001101111000100000111000000;
filter5[9][501] = 35'b11111110111111010101110100110000000;
filter5[9][502] = 35'b11111101111110100101110100011000000;
filter5[9][503] = 35'b00000000100001000110011000111011000;
filter5[9][504] = 35'b11111111000011100110101001011111000;
filter5[9][505] = 35'b00000000100010010110011001000010000;
filter5[9][506] = 35'b11111101111111101000001001100000000;
filter5[9][507] = 35'b00000001001111011101100101101110000;
filter5[9][508] = 35'b00000010111111000010110011111100000;
filter5[9][509] = 35'b00000000011110111110011000000111000;
filter5[9][510] = 35'b11111111000111001110100011011001000;
filter5[9][511] = 35'b11111111101110110010111010010101100;
filter5[9][512] = 35'b00000001000101000110010110100110000;
filter5[9][513] = 35'b00000001011010101010110001010100000;
filter5[9][514] = 35'b11111111101101000011001000110111100;
filter5[9][515] = 35'b11111010010111011111110000010000000;
filter5[9][516] = 35'b11111110101001101010111101101010000;
filter5[9][517] = 35'b11111110100110101000110110101010000;
filter5[9][518] = 35'b00000001010010111011000010101010000;
filter5[9][519] = 35'b00000001100010101111101110101110000;
filter5[9][520] = 35'b00000000001100011111001001110011000;
filter5[9][521] = 35'b11111111110010001101011010101101100;
filter5[9][522] = 35'b00000000010111101111100000101011100;
filter5[9][523] = 35'b00000010101101001011011111000100000;
filter5[9][524] = 35'b00000000111010100001011000001000000;
filter5[9][525] = 35'b11111110111000001010000010010110000;
filter5[9][526] = 35'b11111011111100110010011111100000000;
filter5[9][527] = 35'b00000000101100000101101111001011000;
filter5[9][528] = 35'b00000000000110011010101010000000111;
filter5[9][529] = 35'b11111011001001011100111001010000000;
filter5[9][530] = 35'b00000000010010111100010110100010000;
filter5[9][531] = 35'b00000001010110111001101111010100000;
filter5[9][532] = 35'b00000001011110101111101011111000000;
filter5[9][533] = 35'b11111111010001001010100110100111000;
filter5[9][534] = 35'b11111011111110001101110000001000000;
filter5[9][535] = 35'b11111110110011101111101101100000000;
filter5[9][536] = 35'b00000000000011011101001010010101010;
filter5[9][537] = 35'b11111101110101101001010110011100000;
filter5[9][538] = 35'b11111110010001110010001011110110000;
filter5[9][539] = 35'b00000000111111111001110110100101000;
filter5[9][540] = 35'b11111111111001011110010011100011101;
filter5[9][541] = 35'b11111101011101110101011100100100000;
filter5[9][542] = 35'b00000010100000000010010101000000000;
filter5[9][543] = 35'b11111111100101001010011100000010100;
filter5[9][544] = 35'b00000011110100101100010001100000000;
filter5[9][545] = 35'b11111111001100000111011010111000000;
filter5[9][546] = 35'b00000000000101101111111101001000101;
filter5[9][547] = 35'b11111111110110010011110101101010100;
filter5[9][548] = 35'b00000100010011001101101111000000000;
filter5[9][549] = 35'b00000000001001001100000111010010100;
filter5[9][550] = 35'b00000010011101000101100110101000000;
filter5[9][551] = 35'b11111111011100100000100110001101000;
filter5[9][552] = 35'b11111110011000010101010001011100000;
filter5[9][553] = 35'b00000000001001010000011111111000110;
filter5[9][554] = 35'b00000100110100010110010001011000000;
filter5[9][555] = 35'b00000010110100111110100101110000000;
filter5[9][556] = 35'b00000010100000111111100111101100000;
filter5[9][557] = 35'b11111110101101001000100010100100000;
filter5[9][558] = 35'b00000010001111011101101011100000000;
filter5[9][559] = 35'b11111110101001100000110011101000000;
filter5[9][560] = 35'b00000111000101100111000111010000000;
filter5[9][561] = 35'b11111111000000101001111011011001000;
filter5[9][562] = 35'b11111110111011100110010011011000000;
filter5[9][563] = 35'b00000001011111111110010111001010000;
filter5[9][564] = 35'b11111110101111000011010011110000000;
filter5[9][565] = 35'b11111001011110110100110100100000000;
filter5[9][566] = 35'b00000000111000110100100011001000000;
filter5[9][567] = 35'b00000001110010011110010001011110000;
filter5[9][568] = 35'b11111110101011010001111101110110000;
filter5[9][569] = 35'b00000001101101011001110110111110000;
filter5[9][570] = 35'b11111111011001000011101101000111000;
filter5[9][571] = 35'b11111110100001111111100111001000000;
filter5[9][572] = 35'b11111110100100111100000111010000000;
filter5[9][573] = 35'b11111100000111000101000001101100000;
filter5[9][574] = 35'b11111110111011110011111001100100000;
filter5[9][575] = 35'b00000001101000001011111110001010000;
filter5[9][576] = 35'b00000000101001010001010110101010000;
filter5[9][577] = 35'b00000001000111101010010000100110000;
filter5[9][578] = 35'b00000001101010101100111101101110000;
filter5[9][579] = 35'b11111111001000001011010111011100000;
filter5[9][580] = 35'b11111110100101100001000010110100000;
filter5[9][581] = 35'b11111101111011101001000101100100000;
filter5[9][582] = 35'b00000011100100110011000111011100000;
filter5[9][583] = 35'b11111101011111001101111100111000000;
filter5[9][584] = 35'b11111101000011010011000110110100000;
filter5[9][585] = 35'b00000001111101111101100010010000000;
filter5[9][586] = 35'b00000010010101100110100101000000000;
filter5[9][587] = 35'b11111111101101101111011010011011100;
filter5[9][588] = 35'b00000010000100000100111100011000000;
filter5[9][589] = 35'b11111101101011110111111100001100000;
filter5[9][590] = 35'b11111011100110111111000011100000000;
filter5[9][591] = 35'b00000011101100111100100111010000000;
filter5[9][592] = 35'b00000100000011000110011100111000000;
filter5[9][593] = 35'b00000000011111000011011110010101000;
filter5[9][594] = 35'b11111110100000010100111011001110000;
filter5[9][595] = 35'b00000001111010011101000100110000000;
filter5[9][596] = 35'b00000001000110110010100011100110000;
filter5[9][597] = 35'b11111111100001101111100110011000100;
filter5[9][598] = 35'b11111001110001011011000111010000000;
filter5[9][599] = 35'b11111110101001101100101000100110000;
filter5[9][600] = 35'b11111101001010001011011011010100000;
filter5[9][601] = 35'b00000001100010111010101000110100000;
filter5[9][602] = 35'b11111111010100000011100010101100000;
filter5[9][603] = 35'b11111100010100001011010000100100000;
filter5[9][604] = 35'b11111110111100000000101011100000000;
filter5[9][605] = 35'b11111110101101111000111100100010000;
filter5[9][606] = 35'b11111101010000011001110110001000000;
filter5[9][607] = 35'b00000000011100100111010101111110000;
filter5[9][608] = 35'b11111101011100011011100011011000000;
filter5[9][609] = 35'b00000010101010101110011101001000000;
filter5[9][610] = 35'b11111111000100111010101100110010000;
filter5[9][611] = 35'b11111101101011000110100100011000000;
filter5[9][612] = 35'b00000001000001111101101000101000000;
filter5[9][613] = 35'b11111110101011001000010001011100000;
filter5[9][614] = 35'b00000001111111010001011000111110000;
filter5[9][615] = 35'b00000010000110010010101100100000000;
filter5[9][616] = 35'b00000000010011110110101110000011100;
filter5[9][617] = 35'b00000000010111010011000111010000000;
filter5[9][618] = 35'b00000101010000110100000101010000000;
filter5[9][619] = 35'b00000000100111010001100101110010000;
filter5[9][620] = 35'b00000010100010010100100000101100000;
filter5[9][621] = 35'b11111111101010010011001110111011000;
filter5[9][622] = 35'b00000001001111100101100100110100000;
filter5[9][623] = 35'b00000000111001001100100101001011000;
filter5[9][624] = 35'b00000001110101111101101011011110000;
filter5[9][625] = 35'b11111111001101111011110110111100000;
filter5[9][626] = 35'b11111100110000011011010101111000000;
filter5[9][627] = 35'b11111100000001001001100110011000000;
filter5[9][628] = 35'b00000011101111111110000001101000000;
filter5[9][629] = 35'b11111010100100110101111011011000000;
filter5[9][630] = 35'b11111110101001000000100001110000000;
filter5[9][631] = 35'b00000011000111000110100111100100000;
filter5[9][632] = 35'b00000111000001011000010000010000000;
filter5[9][633] = 35'b00000000010000010000101010011101000;
filter5[9][634] = 35'b11111110101001110101011000110010000;
filter5[9][635] = 35'b00000100101111011010111011111000000;
filter5[9][636] = 35'b00000011010000000100010011001000000;
filter5[9][637] = 35'b11111111101010011001101100111110100;
filter5[9][638] = 35'b00000001010111111010101011101100000;
filter5[9][639] = 35'b11111100101100011110001001101000000;
filter5[9][640] = 35'b11111100010001010010111010111100000;
filter5[9][641] = 35'b11111110011001101101111111011000000;
filter5[9][642] = 35'b11111111101101001001110111010010000;
filter5[9][643] = 35'b00000000000000011110010101010001010;
filter5[9][644] = 35'b11111101000110100010001110000100000;
filter5[9][645] = 35'b00000010010001101100001000010000000;
filter5[9][646] = 35'b00000000100101100100100111100101000;
filter5[9][647] = 35'b11111111101001011101110100100010000;
filter5[9][648] = 35'b00000000011001101011000101001000000;
filter5[9][649] = 35'b00000010110010000000101110111100000;
filter5[9][650] = 35'b11111010111110110101001111100000000;
filter5[9][651] = 35'b00000001100100111010100000000100000;
filter5[9][652] = 35'b00000011110101101000000001011100000;
filter5[9][653] = 35'b00000011011011111110101100101000000;
filter5[9][654] = 35'b11111110001001101010100110101000000;
filter5[9][655] = 35'b00000011110100101101110111110100000;
filter5[9][656] = 35'b11111101101010000000000000100000000;
filter5[9][657] = 35'b11111100010111010000111010010100000;
filter5[9][658] = 35'b11111111001101110100000010111010000;
filter5[9][659] = 35'b00000010000000111111101101011100000;
filter5[9][660] = 35'b11111110101111110101000011110100000;
filter5[9][661] = 35'b11111011110000010101011000100000000;
filter5[9][662] = 35'b00000011111101001100100010101000000;
filter5[9][663] = 35'b11111111110011000110110110100011000;
filter5[9][664] = 35'b00000000100100111111010101010111000;
filter5[9][665] = 35'b11111010000000110110101110000000000;
filter5[9][666] = 35'b11111101000101010100001001011100000;
filter5[9][667] = 35'b11111110011111000011001111010000000;
filter5[9][668] = 35'b00000000001101100010111001110110010;
filter5[9][669] = 35'b11111111101100110101100111011100100;
filter5[9][670] = 35'b11111110011111110111101111101000000;
filter5[9][671] = 35'b00000000100000000010111011101110000;
filter5[9][672] = 35'b11111110101100011101000110011100000;
filter5[9][673] = 35'b00000010000100110111011101011000000;
filter5[9][674] = 35'b00000100000110100111001000011000000;
filter5[9][675] = 35'b11111110100110100101101100000010000;
filter5[9][676] = 35'b00000010001001101011011111010000000;
filter5[9][677] = 35'b11111011100000011010110111000000000;
filter5[9][678] = 35'b00000010010101000100000100111100000;
filter5[9][679] = 35'b11111110001110100100010011110010000;
filter5[9][680] = 35'b11111011010000110110011110010000000;
filter5[9][681] = 35'b11111110000110110111100001111000000;
filter5[9][682] = 35'b00000101101111001101000100011000000;
filter5[9][683] = 35'b00000000101000010101010000111100000;
filter5[9][684] = 35'b11111110100100001011101110100000000;
filter5[9][685] = 35'b00000000001100101011001111100110110;
filter5[9][686] = 35'b00000001010010101110011010000100000;
filter5[9][687] = 35'b00000101001100001110010111100000000;
filter5[9][688] = 35'b00001000000110010000010111000000000;
filter5[9][689] = 35'b11111111000101000010001111100110000;
filter5[9][690] = 35'b00000011100111101111010000011100000;
filter5[9][691] = 35'b00000000101100101110010111110100000;
filter5[9][692] = 35'b00000010101100011111111010001000000;
filter5[9][693] = 35'b11111100010101001011101110100100000;
filter5[9][694] = 35'b11111111101100010000000001011000100;
filter5[9][695] = 35'b11111100001011110110100100111100000;
filter5[9][696] = 35'b11111111110011101100000111100001000;
filter5[9][697] = 35'b00000001110101100100010000010010000;
filter5[9][698] = 35'b11111111111111011110011110010010100;
filter5[9][699] = 35'b11111110001111010101101010001010000;
filter5[9][700] = 35'b11111110000001100001111101100100000;
filter5[9][701] = 35'b00000010101010010000110111010000000;
filter5[9][702] = 35'b00000010011010110111001001100100000;
filter5[9][703] = 35'b00000001110000011011100001001110000;
filter5[9][704] = 35'b11111101100101000111011100111100000;
filter5[9][705] = 35'b11111111101110111001110111001100100;
filter5[9][706] = 35'b00000000011100010111010101011000000;
filter5[9][707] = 35'b11111111010000110001111001010010000;
filter5[9][708] = 35'b11111111100010110000110010000101100;
filter5[9][709] = 35'b11111111001110011110100101100011000;
filter5[9][710] = 35'b11111111100110000010100110111101000;
filter5[9][711] = 35'b11111110101100101001001110001010000;
filter5[9][712] = 35'b11111111100001100100100001001110100;
filter5[9][713] = 35'b11111111101111011100010111011111100;
filter5[9][714] = 35'b00000000110001011111000011000000000;
filter5[9][715] = 35'b11111110011001000100101000010000000;
filter5[9][716] = 35'b11111110011110101110110101001100000;
filter5[9][717] = 35'b00000000011100011000101000110000000;
filter5[9][718] = 35'b00000000011101111000000001010110000;
filter5[9][719] = 35'b00000001000001010111001100101110000;
filter5[9][720] = 35'b11111110110111000110010100100110000;
filter5[9][721] = 35'b11111111111100011010010100101111100;
filter5[9][722] = 35'b11111101111111011110111100010100000;
filter5[9][723] = 35'b00000000100001111110100100110111000;
filter5[9][724] = 35'b00000011101011100110100011110000000;
filter5[9][725] = 35'b11111100000111111000110101011000000;
filter5[9][726] = 35'b11111111011000000100101010000010000;
filter5[9][727] = 35'b11111110101100010001011111010110000;
filter5[9][728] = 35'b00000000001110001111100001001111110;
filter5[9][729] = 35'b11111101001011000001111001010000000;
filter5[9][730] = 35'b11111101111001110111011001000000000;
filter5[9][731] = 35'b11111110111000010111100100101110000;
filter5[9][732] = 35'b00000000011010111011110101000010000;
filter5[9][733] = 35'b11111110100011000001011101000010000;
filter5[9][734] = 35'b11111100001010010001010110110100000;
filter5[9][735] = 35'b11111011111001100111101010100000000;
filter5[9][736] = 35'b00000000010001101101101101111110100;
filter5[9][737] = 35'b11111011001000010011111010101000000;
filter5[9][738] = 35'b11111101100001001011011010000000000;
filter5[9][739] = 35'b11111101010011100000000111001100000;
filter5[9][740] = 35'b00000001110011000100001011000010000;
filter5[9][741] = 35'b11111100110001110100000110001000000;
filter5[9][742] = 35'b11111110100010000000100010110000000;
filter5[9][743] = 35'b00000010100001000111101100010100000;
filter5[9][744] = 35'b00000101011101010101100111101000000;
filter5[9][745] = 35'b11111101100000010111011000010100000;
filter5[9][746] = 35'b11111110011010111011111100101000000;
filter5[9][747] = 35'b11111101010011110011001010111100000;
filter5[9][748] = 35'b11111110101011001011010000111000000;
filter5[9][749] = 35'b11111101100011010101110111011000000;
filter5[9][750] = 35'b00001000101011111000001000110000000;
filter5[9][751] = 35'b00000000111000100001011011010001000;
filter5[9][752] = 35'b00000000011110101011100001110110100;
filter5[9][753] = 35'b00000000101010111100101111011000000;
filter5[9][754] = 35'b00000011011001011011000111100100000;
filter5[9][755] = 35'b00000100001110100010010011101000000;
filter5[9][756] = 35'b00000010010010011110000000010000000;
filter5[9][757] = 35'b11111110000011111110100111010100000;
filter5[9][758] = 35'b00000011100001110101011110011000000;
filter5[9][759] = 35'b11111111001111110000110001001010000;
filter5[9][760] = 35'b11111100111000100100001101101000000;
filter5[9][761] = 35'b11111010110011100010011000100000000;
filter5[9][762] = 35'b11111110100110010100110110111010000;
filter5[9][763] = 35'b00000001111101110000000100101010000;
filter5[9][764] = 35'b11111111101010001100010100000011100;
filter5[9][765] = 35'b11111110011101111000111011111010000;
filter5[9][766] = 35'b11111001110010001111000001011000000;
filter5[9][767] = 35'b11111111100001000100101110010001100;
filter5[9][768] = 35'b00000010100100101011111101010100000;
filter5[9][769] = 35'b11111110101111100110100001110110000;
filter5[9][770] = 35'b00000001100011001111000100010100000;
filter5[9][771] = 35'b00000001000011111101011010010010000;
filter5[9][772] = 35'b11111111000000001101011000001100000;
filter5[9][773] = 35'b11111101001111011110010111001000000;
filter5[9][774] = 35'b11111110001100111011010100100100000;
filter5[9][775] = 35'b11111101011011000011010111110100000;
filter5[9][776] = 35'b11111101010011001011001001111000000;
filter5[9][777] = 35'b00000000000101011110000101011100011;
filter5[9][778] = 35'b11111111000111000111110111110111000;
filter5[9][779] = 35'b00000010011111110110011100000100000;
filter5[9][780] = 35'b11111110000000111111000000001110000;
filter5[9][781] = 35'b11111110000000010100011110101000000;
filter5[9][782] = 35'b00000001101111111000111100001100000;
filter5[9][783] = 35'b11111111000001000000111101010110000;
filter5[9][784] = 35'b11111101110000010110100110000100000;
filter5[9][785] = 35'b11111110101101001010001100101100000;
filter5[9][786] = 35'b00000001101010011011010010111100000;
filter5[9][787] = 35'b11111011101110010101000111000000000;
filter5[9][788] = 35'b00000100001111110001111011110000000;
filter5[9][789] = 35'b00000010111000100100010011110100000;
filter5[9][790] = 35'b00000001001100000001100101111110000;
filter5[9][791] = 35'b11111100110011010110011101010000000;
filter5[9][792] = 35'b11111100000110000111111111000100000;
filter5[9][793] = 35'b00000000011101001100100001000000000;
filter5[9][794] = 35'b11111011111111000101110010000000000;
filter5[9][795] = 35'b11111111100010001110111001100000100;
filter5[9][796] = 35'b11111001000100001110110100111000000;
filter5[9][797] = 35'b11111111111111101101011101100111010;
filter5[9][798] = 35'b00001000011000101101001011010000000;
filter5[9][799] = 35'b11110100010000011001000100110000000;
filter5[9][800] = 35'b00000000100010001001111110000010000;
filter5[9][801] = 35'b00000001010010001110100001111100000;
filter5[9][802] = 35'b11111010111100100100111110111000000;
filter5[9][803] = 35'b11111001101001101011111000011000000;
filter5[9][804] = 35'b00000000110111110111011101101001000;
filter5[9][805] = 35'b00000011000011011111101100011100000;
filter5[9][806] = 35'b00000111011110101110010101010000000;
filter5[9][807] = 35'b00000111011100101110111010101000000;
filter5[9][808] = 35'b11111101111010110100001000000000000;
filter5[9][809] = 35'b00000010001001111111111010111000000;
filter5[9][810] = 35'b00000000010001000001010001001101100;
filter5[9][811] = 35'b00000011111011111100110110001000000;
filter5[9][812] = 35'b11111101010110010010010010101000000;
filter5[9][813] = 35'b00001010101001101110101010100000000;
filter5[9][814] = 35'b00000010111101010010101101111100000;
filter5[9][815] = 35'b11111110000100101111110100010100000;
filter5[9][816] = 35'b00000000101010110111101100001001000;
filter5[9][817] = 35'b00000010110001010000101110011100000;
filter5[9][818] = 35'b11111000001110100111011001111000000;
filter5[9][819] = 35'b11111111100110101100110101010111000;
filter5[9][820] = 35'b00000110011100011000010100000000000;
filter5[9][821] = 35'b00000000011110010110000011000100000;
filter5[9][822] = 35'b00000010001011011001001110101100000;
filter5[9][823] = 35'b00000010111110111111001011100000000;
filter5[9][824] = 35'b00000011000001011000100101110000000;
filter5[9][825] = 35'b11111101110000001010010100110100000;
filter5[9][826] = 35'b11111110110100111111001000010010000;
filter5[9][827] = 35'b11111110111011110110100111000110000;
filter5[9][828] = 35'b00000000001100001100011111110001000;
filter5[9][829] = 35'b00000000000001101101111000001111001;
filter5[9][830] = 35'b11111110101011011110111111011100000;
filter5[9][831] = 35'b11111011001111111011100110100000000;
filter5[9][832] = 35'b11111101010001000101001000101100000;
filter5[9][833] = 35'b11111111000010001111111101111000000;
filter5[9][834] = 35'b11111110111001110011001000110000000;
filter5[9][835] = 35'b11111110101001011100111101111110000;
filter5[9][836] = 35'b11111101100111111100010101101000000;
filter5[9][837] = 35'b11111111100111101000001111110011100;
filter5[9][838] = 35'b00000000011111101101011101111111100;
filter5[9][839] = 35'b11111111000000011110110101010100000;
filter5[9][840] = 35'b11111111111110101101000101101010011;
filter5[9][841] = 35'b00000000011011011011011010010010000;
filter5[9][842] = 35'b11111110110010010100000000001100000;
filter5[9][843] = 35'b00000000100010011100111111110010000;
filter5[9][844] = 35'b11111111110001101001101010010110110;
filter5[9][845] = 35'b00000000100111011010000111111101000;
filter5[9][846] = 35'b00000000001100011100011000011111100;
filter5[9][847] = 35'b00000000011011011110100101111100000;
filter5[9][848] = 35'b11111111011011100110011001001000000;
filter5[9][849] = 35'b11111111000000110001001010100101000;
filter5[9][850] = 35'b11111111110000100001110101000000000;
filter5[9][851] = 35'b11111110100101111111100010101000000;
filter5[9][852] = 35'b11111011110000011000000111101000000;
filter5[9][853] = 35'b11111110001000101001001010111110000;
filter5[9][854] = 35'b11111111111100000011010111111101011;
filter5[9][855] = 35'b00000000010111011011001111010000100;
filter5[9][856] = 35'b00000000101000000011000010110000000;
filter5[9][857] = 35'b11111101111100101101011010110000000;
filter5[9][858] = 35'b11111110101111001010011101111010000;
filter5[9][859] = 35'b00000000111000011101010011000000000;
filter5[9][860] = 35'b00000101001110011011000110101000000;
filter5[9][861] = 35'b11111111011001101100101000010000000;
filter5[9][862] = 35'b11111100101011101100101100111000000;
filter5[9][863] = 35'b11111111000111101011001110011110000;
filter5[9][864] = 35'b11111111101110010010101001111000000;
filter5[9][865] = 35'b11111110001011101010100000000110000;
filter5[9][866] = 35'b11111100111011101111001000101000000;
filter5[9][867] = 35'b11111111110011111110010101010110100;
filter5[9][868] = 35'b11111101101000010110101101010000000;
filter5[9][869] = 35'b11111100111101100000111001000000000;
filter5[9][870] = 35'b00000000100010010010001110011110000;
filter5[9][871] = 35'b11111101101010111101001000111000000;
filter5[9][872] = 35'b00000001111010110111000100011110000;
filter5[9][873] = 35'b11111110110110011111101001101010000;
filter5[9][874] = 35'b11111100000111100011101110101100000;
filter5[9][875] = 35'b11111110100110101010001011101010000;
filter5[9][876] = 35'b11111111110100011010001001010111110;
filter5[9][877] = 35'b11111110110110100101100100011000000;
filter5[9][878] = 35'b00000100000010011100101000011000000;
filter5[9][879] = 35'b00000100010110001000011111100000000;
filter5[9][880] = 35'b11111110000111010001000111001000000;
filter5[9][881] = 35'b00000001100000000111100010100100000;
filter5[9][882] = 35'b00000011100111101100110111000000000;
filter5[9][883] = 35'b00000001110010000111101001111000000;
filter5[9][884] = 35'b11111111010110011011000101110001000;
filter5[9][885] = 35'b11111101011110100000111010100000000;
filter5[9][886] = 35'b11111110011100010100100100010100000;
filter5[9][887] = 35'b00000000000010000111110001001111101;
filter5[9][888] = 35'b11111010110011110000001000110000000;
filter5[9][889] = 35'b00000000110101000110111000001111000;
filter5[9][890] = 35'b11111101010001011000110111101100000;
filter5[9][891] = 35'b00000111110000111011011100111000000;
filter5[9][892] = 35'b00000001001010011101111100101100000;
filter5[9][893] = 35'b11111001001100110000110000001000000;
filter5[9][894] = 35'b11111101000000111111001011101100000;
filter5[9][895] = 35'b11111101010110100011100000010100000;
filter5[9][896] = 35'b11111101111100100011111011111000000;
filter5[9][897] = 35'b11111000100110111001011101000000000;
filter5[9][898] = 35'b11111010101110010000000110110000000;
filter5[9][899] = 35'b11111010010100111011000010110000000;
filter5[9][900] = 35'b11111101011101111001001011101000000;
filter5[9][901] = 35'b11111100111001101101011100001000000;
filter5[9][902] = 35'b00000000010001101010111011011111100;
filter5[9][903] = 35'b11111011000011010001111011110000000;
filter5[9][904] = 35'b11111011101100010001000000111000000;
filter5[9][905] = 35'b00000001011111010100111111111110000;
filter5[9][906] = 35'b11111010111111100000101001100000000;
filter5[9][907] = 35'b11111100101010111101111111110000000;
filter5[9][908] = 35'b11111001000001000010001011101000000;
filter5[9][909] = 35'b11111101001111111010110000110100000;
filter5[9][910] = 35'b11111001010011110001000010100000000;
filter5[9][911] = 35'b11111101001000110110010010011100000;
filter5[9][912] = 35'b11111100111010100101110011100100000;
filter5[9][913] = 35'b11111000111010101010111100110000000;
filter5[9][914] = 35'b11111011101001000101100100011000000;
filter5[9][915] = 35'b11111100101011110110110000011000000;
filter5[9][916] = 35'b11111110010101001110111010100110000;
filter5[9][917] = 35'b11111010011110110010000111100000000;
filter5[9][918] = 35'b00000010000000100010011011010000000;
filter5[9][919] = 35'b11110111011110001010101011010000000;
filter5[9][920] = 35'b00000111111000001101100101000000000;
filter5[9][921] = 35'b11111101010010001011110010100100000;
filter5[9][922] = 35'b11111100100101101000100011100000000;
filter5[9][923] = 35'b11111111011001111111001111101100000;
filter5[9][924] = 35'b00000111101101100100011000000000000;
filter5[9][925] = 35'b11111010111110100110001111110000000;
filter5[9][926] = 35'b11111111010101000011000110100011000;
filter5[9][927] = 35'b11110000001111001101100100110000000;
filter5[9][928] = 35'b00000010011110001010110000011000000;
filter5[9][929] = 35'b11111000011111010101001011011000000;
filter5[9][930] = 35'b11111011111000001100010110101000000;
filter5[9][931] = 35'b11111101001010010100001000000100000;
filter5[9][932] = 35'b11111111101101101001111000001110000;
filter5[9][933] = 35'b11111100110101100101110110100100000;
filter5[9][934] = 35'b11111110111001100000110011110000000;
filter5[9][935] = 35'b00001010001110010111111001100000000;
filter5[9][936] = 35'b00000111010001100001100111111000000;
filter5[9][937] = 35'b00000001000010111011010100110010000;
filter5[9][938] = 35'b00000001111001010010111101010100000;
filter5[9][939] = 35'b11111011100111100000111010001000000;
filter5[9][940] = 35'b00000000110011011000100110011100000;
filter5[9][941] = 35'b00000000110001011010101111001111000;
filter5[9][942] = 35'b00000001101010000100011100000000000;
filter5[9][943] = 35'b11111111010001110001010000111001000;
filter5[9][944] = 35'b11111110100010111110111000100100000;
filter5[9][945] = 35'b11111101011011001110110111110100000;
filter5[9][946] = 35'b00000001000101011111001100100000000;
filter5[9][947] = 35'b00000100000010001010000111001000000;
filter5[9][948] = 35'b11111100011111011101111001001000000;
filter5[9][949] = 35'b11111110110000101001000011110110000;
filter5[9][950] = 35'b11111011100001100100110011110000000;
filter5[9][951] = 35'b11111011011010001010011100000000000;
filter5[9][952] = 35'b11111011110111000010001101000000000;
filter5[9][953] = 35'b11111101010110110000010101011000000;
filter5[9][954] = 35'b00000010100010100101101101000100000;
filter5[9][955] = 35'b00000100011010101101000101000000000;
filter5[9][956] = 35'b00000010010001010001000000000000000;
filter5[9][957] = 35'b11111011010011110010011111111000000;
filter5[9][958] = 35'b11101011111111001101010111000000000;
filter5[9][959] = 35'b11111100000010110011010001101100000;
filter5[9][960] = 35'b00000011101000010011110011011000000;
filter5[9][961] = 35'b11111110111010011001110110100000000;
filter5[9][962] = 35'b00000001010000110110111110000010000;
filter5[9][963] = 35'b00000000111011111001010001000100000;
filter5[9][964] = 35'b11111000110100101000100011001000000;
filter5[9][965] = 35'b00000011000100001000101111011100000;
filter5[9][966] = 35'b00000101010011001110011100000000000;
filter5[9][967] = 35'b00000100111110110101100010010000000;
filter5[9][968] = 35'b00000000110110011011101001111100000;
filter5[9][969] = 35'b00000000011101001010110101010001100;
filter5[9][970] = 35'b11111111110010110101001010110010100;
filter5[9][971] = 35'b11111100110110111001010010110000000;
filter5[9][972] = 35'b11111011001000100011100111111000000;
filter5[9][973] = 35'b11111110011111011111001101001000000;
filter5[9][974] = 35'b11111100101011100001110100010100000;
filter5[9][975] = 35'b00000011100001010000111001100000000;
filter5[9][976] = 35'b00000000101100001110100111110010000;
filter5[9][977] = 35'b11111101110011110100000000011100000;
filter5[9][978] = 35'b11101110110000010010100100100000000;
filter5[9][979] = 35'b00000011011101010111100111000000000;
filter5[9][980] = 35'b00000010011101001110000010111100000;
filter5[9][981] = 35'b00000000000001110001100010110001000;
filter5[9][982] = 35'b00000100000111011000110110101000000;
filter5[9][983] = 35'b00000001010000001001100110110110000;
filter5[9][984] = 35'b00001000110000101101101010100000000;
filter5[9][985] = 35'b00000111000111110010011010000000000;
filter5[9][986] = 35'b11111011000000111100111000111000000;
filter5[9][987] = 35'b11111111110011110010111100111010010;
filter5[9][988] = 35'b00000010110001111110100000001100000;
filter5[9][989] = 35'b00000001000010010010011001011000000;
filter5[9][990] = 35'b11111111110000001001001101110110100;
filter5[9][991] = 35'b00000000100111010100110111101110000;
filter5[9][992] = 35'b00000100010010111011010110101000000;
filter5[9][993] = 35'b11111101011101111111100000001100000;
filter5[9][994] = 35'b11111010001010110110110000100000000;
filter5[9][995] = 35'b11111101011110111111000101000100000;
filter5[9][996] = 35'b00000001010100101010010001101100000;
filter5[9][997] = 35'b11111011101010100100000010000000000;
filter5[9][998] = 35'b11111111111101001101111110000010111;
filter5[9][999] = 35'b00000001111011100000000001110000000;
filter5[9][1000] = 35'b00001010110101111111101000100000000;
filter5[9][1001] = 35'b00000110001100100010010011010000000;
filter5[9][1002] = 35'b00000001000101100101100100101010000;
filter5[9][1003] = 35'b11111110001110110101001111000010000;
filter5[9][1004] = 35'b00000001100110110001101110010100000;
filter5[9][1005] = 35'b11111100110000010100010110000000000;
filter5[9][1006] = 35'b11111111100011111110011101000011100;
filter5[9][1007] = 35'b00000011000110100010101110110000000;
filter5[9][1008] = 35'b11111011111110001101010110110000000;
filter5[9][1009] = 35'b11111011110010000001100111011000000;
filter5[9][1010] = 35'b11111101011001011111110110111000000;
filter5[9][1011] = 35'b00000011010001111110101010111100000;
filter5[9][1012] = 35'b11111110111010000101010010001000000;
filter5[9][1013] = 35'b11110100001011011111111100110000000;
filter5[9][1014] = 35'b00000110100000000011010001110000000;
filter5[9][1015] = 35'b00000011111101001111111111011100000;
filter5[9][1016] = 35'b00000000010100110011100000011101000;
filter5[9][1017] = 35'b11111110011110011110110010011000000;
filter5[9][1018] = 35'b00000101010100110010001101000000000;
filter5[9][1019] = 35'b00000111001001000111100110000000000;
filter5[9][1020] = 35'b11111110100000011110011100011000000;
filter5[9][1021] = 35'b11111000111011001100110101100000000;
filter5[9][1022] = 35'b11110101010110101110100010000000000;
filter5[9][1023] = 35'b11111100110010110110111010011100000;
filter5[10][0] = 35'b11111010010001001001100010100000000;
filter5[10][1] = 35'b00000100101000010101011011000000000;
filter5[10][2] = 35'b00000001110100011101110001101110000;
filter5[10][3] = 35'b00000100000001101000001100001000000;
filter5[10][4] = 35'b11111100111001011001110100111000000;
filter5[10][5] = 35'b00000001010100101101111100001000000;
filter5[10][6] = 35'b00000110011010101010011111011000000;
filter5[10][7] = 35'b11111110011110110000111110011010000;
filter5[10][8] = 35'b00000100000000000101010000101000000;
filter5[10][9] = 35'b11111101101100111001110011000000000;
filter5[10][10] = 35'b00000000101011111110110010110001000;
filter5[10][11] = 35'b11111100111111011101001011111100000;
filter5[10][12] = 35'b11111100111010011101001101100000000;
filter5[10][13] = 35'b11111101111111010010101111001000000;
filter5[10][14] = 35'b00000001010101111110110000011010000;
filter5[10][15] = 35'b11111000100001111011001111100000000;
filter5[10][16] = 35'b00000000010110101001000000000011000;
filter5[10][17] = 35'b11111100100010001111101101111000000;
filter5[10][18] = 35'b11111110110101011111001011110100000;
filter5[10][19] = 35'b00000010011101110110101000101000000;
filter5[10][20] = 35'b11111111011011001101011101110011000;
filter5[10][21] = 35'b00000001001001001110111000011010000;
filter5[10][22] = 35'b11111010011010011111000111001000000;
filter5[10][23] = 35'b11111000101011111010111101111000000;
filter5[10][24] = 35'b11111110110100001000110101101100000;
filter5[10][25] = 35'b11111111010010010000110110100001000;
filter5[10][26] = 35'b11111110111000001100001011011100000;
filter5[10][27] = 35'b11111100111001011000101000001000000;
filter5[10][28] = 35'b11111110100000101001110011000100000;
filter5[10][29] = 35'b00000101100111100111010001011000000;
filter5[10][30] = 35'b11111110001110010110011110110000000;
filter5[10][31] = 35'b00000100011010001001100110100000000;
filter5[10][32] = 35'b00000000011010010100101001100100000;
filter5[10][33] = 35'b00000000100111101011000001010100000;
filter5[10][34] = 35'b00000001000001100101111111111010000;
filter5[10][35] = 35'b11111111010011001101001111010001000;
filter5[10][36] = 35'b11111100100111011010101100111100000;
filter5[10][37] = 35'b11111110111101000011011110100010000;
filter5[10][38] = 35'b11111001011011011100111011000000000;
filter5[10][39] = 35'b11111101011111001011001001011000000;
filter5[10][40] = 35'b11111110001100111101010101101110000;
filter5[10][41] = 35'b00000000000001000101100110100100011;
filter5[10][42] = 35'b11111110100110110011011001101000000;
filter5[10][43] = 35'b11111111110011000100110010100100010;
filter5[10][44] = 35'b11111100110100111000000100000100000;
filter5[10][45] = 35'b00000010010110010110000011110000000;
filter5[10][46] = 35'b00000010011001111001101010011000000;
filter5[10][47] = 35'b11111011010000111001000001110000000;
filter5[10][48] = 35'b00000010101000100010110000011000000;
filter5[10][49] = 35'b11111111010011100000011000100100000;
filter5[10][50] = 35'b11111110110011100100010011111010000;
filter5[10][51] = 35'b11111111110110011110001110111011100;
filter5[10][52] = 35'b00000110111100101100100100100000000;
filter5[10][53] = 35'b00000001001010001010100001000010000;
filter5[10][54] = 35'b00000111110111000110001101010000000;
filter5[10][55] = 35'b11111111001011000010111100010101000;
filter5[10][56] = 35'b11111000001111000111010000101000000;
filter5[10][57] = 35'b00000111001101111100100010001000000;
filter5[10][58] = 35'b00000000110111011010110010101010000;
filter5[10][59] = 35'b00000100010000100111100101110000000;
filter5[10][60] = 35'b00000010111010100011111000011100000;
filter5[10][61] = 35'b11111111000111001011011110011011000;
filter5[10][62] = 35'b11111011011000111010111011101000000;
filter5[10][63] = 35'b00001100000011101100010110010000000;
filter5[10][64] = 35'b00000010110010110101011001111100000;
filter5[10][65] = 35'b00000111011101010111000001110000000;
filter5[10][66] = 35'b00000101011111000111100100000000000;
filter5[10][67] = 35'b00000100001010001010011101111000000;
filter5[10][68] = 35'b11111100100110101100010011100000000;
filter5[10][69] = 35'b00000010110101111111111001000100000;
filter5[10][70] = 35'b00000010110100000000100010100000000;
filter5[10][71] = 35'b11111110011101111100110011110000000;
filter5[10][72] = 35'b00001010100000110011110001000000000;
filter5[10][73] = 35'b11111111100000001101000111011101100;
filter5[10][74] = 35'b00000000100001000100100110110000000;
filter5[10][75] = 35'b11111110010100000111101011100000000;
filter5[10][76] = 35'b11111110001110110000010001100110000;
filter5[10][77] = 35'b00000001110101111001101110110110000;
filter5[10][78] = 35'b11111111100011011110000000100001000;
filter5[10][79] = 35'b11111100100110011000010001011100000;
filter5[10][80] = 35'b00000001100101111101100111000100000;
filter5[10][81] = 35'b00000000110000110000101101011011000;
filter5[10][82] = 35'b11111101101100110001110110011100000;
filter5[10][83] = 35'b11111111011101110001000110111110000;
filter5[10][84] = 35'b00000000000000001111100011101011110;
filter5[10][85] = 35'b00000000010111001011100100010111100;
filter5[10][86] = 35'b00000001010001100101101101100010000;
filter5[10][87] = 35'b11111000011101111100001000101000000;
filter5[10][88] = 35'b11111111000010010011100011111011000;
filter5[10][89] = 35'b00000001101111010010000000100110000;
filter5[10][90] = 35'b11111100101011110100000010001000000;
filter5[10][91] = 35'b11111011001110000110001110000000000;
filter5[10][92] = 35'b00000100001001100001101010000000000;
filter5[10][93] = 35'b00000010111111000110001011110000000;
filter5[10][94] = 35'b11111101100000011000100011011100000;
filter5[10][95] = 35'b00000100001101101011011001001000000;
filter5[10][96] = 35'b11111111111111110100101101100010101;
filter5[10][97] = 35'b00000000101101000111101011010010000;
filter5[10][98] = 35'b00000000111101100000000111100011000;
filter5[10][99] = 35'b11111001111100100100000001001000000;
filter5[10][100] = 35'b11111101111111100100000110111000000;
filter5[10][101] = 35'b11111110000011100000101011010110000;
filter5[10][102] = 35'b11111101010101111100011100100000000;
filter5[10][103] = 35'b00000100101110010100011001011000000;
filter5[10][104] = 35'b00000000001100101010111110100111010;
filter5[10][105] = 35'b00000010111101000100110010100000000;
filter5[10][106] = 35'b11111111011010111001001000010001000;
filter5[10][107] = 35'b00000001100011100100011011101010000;
filter5[10][108] = 35'b11111111000000000100001100010110000;
filter5[10][109] = 35'b00000010000000000011100010000100000;
filter5[10][110] = 35'b11111101000011101000011111101000000;
filter5[10][111] = 35'b11111101011111000100100001111000000;
filter5[10][112] = 35'b00000011110001001010111011111100000;
filter5[10][113] = 35'b11111110110010001001010110101100000;
filter5[10][114] = 35'b11111111001110001110100101010000000;
filter5[10][115] = 35'b00000001111110011111001001011000000;
filter5[10][116] = 35'b11111110001001010000000111100010000;
filter5[10][117] = 35'b11111101111000111010000111111000000;
filter5[10][118] = 35'b11111110010100011111100000101100000;
filter5[10][119] = 35'b00000001111111000000100010110110000;
filter5[10][120] = 35'b11111111010011000110011110010001000;
filter5[10][121] = 35'b00000100011100101101101000110000000;
filter5[10][122] = 35'b11111111010100110011001111101111000;
filter5[10][123] = 35'b00000010111101001111001110010000000;
filter5[10][124] = 35'b00000111001001101000011101001000000;
filter5[10][125] = 35'b00000001101111110101110001001010000;
filter5[10][126] = 35'b00000100100110110100111000100000000;
filter5[10][127] = 35'b00001111100100001000101101000000000;
filter5[10][128] = 35'b00010011010111110110110101100000000;
filter5[10][129] = 35'b00001110101000110000010010000000000;
filter5[10][130] = 35'b00000110100001000000111111101000000;
filter5[10][131] = 35'b11111111100000100110111110111111000;
filter5[10][132] = 35'b11111010000101100100010001101000000;
filter5[10][133] = 35'b11111011000111001111110000100000000;
filter5[10][134] = 35'b11111101000010101101111001101100000;
filter5[10][135] = 35'b11110101101000001011010101100000000;
filter5[10][136] = 35'b00010000000100111010000100100000000;
filter5[10][137] = 35'b11111111001001000110111111000100000;
filter5[10][138] = 35'b11111101001011111110100010011000000;
filter5[10][139] = 35'b11111100001001100010000000101100000;
filter5[10][140] = 35'b11111111010001000111111000001001000;
filter5[10][141] = 35'b00000010111100000100111101111000000;
filter5[10][142] = 35'b11111101001000001010011101110100000;
filter5[10][143] = 35'b00000000111000110001010010100010000;
filter5[10][144] = 35'b00000010101101001010110011011000000;
filter5[10][145] = 35'b00000000100110011011111110111110000;
filter5[10][146] = 35'b11111010001000000000011100101000000;
filter5[10][147] = 35'b00000001000110010100101001110000000;
filter5[10][148] = 35'b11111111011000100001110101000010000;
filter5[10][149] = 35'b00000001011101110110101111010110000;
filter5[10][150] = 35'b11111110101110101011110100001010000;
filter5[10][151] = 35'b11111101010010110001011011011000000;
filter5[10][152] = 35'b11111100101100111110001101011100000;
filter5[10][153] = 35'b11111101100010101101011011110100000;
filter5[10][154] = 35'b00000010000010111110111111000100000;
filter5[10][155] = 35'b00000010001001001010000001001000000;
filter5[10][156] = 35'b11111101010000100011010000111100000;
filter5[10][157] = 35'b11111010001010011110000101110000000;
filter5[10][158] = 35'b00000000110010000110010010011111000;
filter5[10][159] = 35'b00001001100011100111101000000000000;
filter5[10][160] = 35'b00000010100100001010100010011000000;
filter5[10][161] = 35'b11111011001000000110100110110000000;
filter5[10][162] = 35'b00000100110011001100101110000000000;
filter5[10][163] = 35'b11111010010111010100110000010000000;
filter5[10][164] = 35'b11111001011000111010100111000000000;
filter5[10][165] = 35'b00000000000100101000000001101111110;
filter5[10][166] = 35'b00000001100000101000110111110100000;
filter5[10][167] = 35'b00000000000110110100000111000000100;
filter5[10][168] = 35'b00000010110011101000110100010000000;
filter5[10][169] = 35'b00000011010100110011000000011000000;
filter5[10][170] = 35'b11111101001100111100010111101000000;
filter5[10][171] = 35'b11111001010101000100000010111000000;
filter5[10][172] = 35'b11111000010000110110101011000000000;
filter5[10][173] = 35'b00000110000010110111110100011000000;
filter5[10][174] = 35'b11111111001000010010100100111101000;
filter5[10][175] = 35'b00001111011101011110000100100000000;
filter5[10][176] = 35'b00010001111011100000000110000000000;
filter5[10][177] = 35'b00000101110100001111000011101000000;
filter5[10][178] = 35'b11110101000110000110010111110000000;
filter5[10][179] = 35'b00000010010110001000011010010000000;
filter5[10][180] = 35'b11111101001010100100011011111100000;
filter5[10][181] = 35'b00000110010010111000011010001000000;
filter5[10][182] = 35'b00000100100110110010001111101000000;
filter5[10][183] = 35'b11111101101011101100001110110000000;
filter5[10][184] = 35'b11110011011000110011111100110000000;
filter5[10][185] = 35'b11111001100010000111010010101000000;
filter5[10][186] = 35'b00010000011010001010110010000000000;
filter5[10][187] = 35'b00000111011000000010011100000000000;
filter5[10][188] = 35'b00001000000110110011100010010000000;
filter5[10][189] = 35'b00011011010101010001010101000000000;
filter5[10][190] = 35'b00000111000101010011100001000000000;
filter5[10][191] = 35'b00001111011100101100001011010000000;
filter5[10][192] = 35'b00000111011101010010011110000000000;
filter5[10][193] = 35'b00000110111100010011011110100000000;
filter5[10][194] = 35'b00001101011110100010010000110000000;
filter5[10][195] = 35'b00000100111011000011011101110000000;
filter5[10][196] = 35'b11101111101001101011100010100000000;
filter5[10][197] = 35'b00000000110100111111110001001011000;
filter5[10][198] = 35'b11111011100010010000011001110000000;
filter5[10][199] = 35'b11110000101011010000001000100000000;
filter5[10][200] = 35'b00000111100001000011001011001000000;
filter5[10][201] = 35'b00001100001100111111011000010000000;
filter5[10][202] = 35'b00000001100101100100000000100100000;
filter5[10][203] = 35'b00000000101000101110011101001011000;
filter5[10][204] = 35'b11111000000000100001110111101000000;
filter5[10][205] = 35'b11111111011100000101001111001100000;
filter5[10][206] = 35'b11111101001111101011010011111100000;
filter5[10][207] = 35'b11111011000101010100000111110000000;
filter5[10][208] = 35'b00000100111101000011101100100000000;
filter5[10][209] = 35'b11111110100100011001001110000100000;
filter5[10][210] = 35'b00000010110101001100010101000000000;
filter5[10][211] = 35'b11111111110101100010101011000000100;
filter5[10][212] = 35'b00000010010101110000110010010000000;
filter5[10][213] = 35'b00000001001011101100001001000000000;
filter5[10][214] = 35'b11111111000101001000001111001001000;
filter5[10][215] = 35'b11111111010001111100011011010000000;
filter5[10][216] = 35'b11111111000100010011111011001101000;
filter5[10][217] = 35'b11111001011000000111011111010000000;
filter5[10][218] = 35'b11111110100110111001110111110100000;
filter5[10][219] = 35'b11111101001011101110101100100000000;
filter5[10][220] = 35'b00000010000010101011011000001000000;
filter5[10][221] = 35'b11111110111011110101110101000110000;
filter5[10][222] = 35'b11111111000111110001110110110010000;
filter5[10][223] = 35'b11111100101101010111011000011100000;
filter5[10][224] = 35'b00000101000101100011101101000000000;
filter5[10][225] = 35'b00000010001110111110100001111100000;
filter5[10][226] = 35'b00000000100101101001101111100000000;
filter5[10][227] = 35'b11111110000110001110010110000000000;
filter5[10][228] = 35'b00000000111000000100100000010110000;
filter5[10][229] = 35'b11111100010001110101110001110100000;
filter5[10][230] = 35'b00000011101110000010110110111100000;
filter5[10][231] = 35'b00000000001100111010101110001001000;
filter5[10][232] = 35'b11110111100011001100000011110000000;
filter5[10][233] = 35'b00000000001100100000001100110000110;
filter5[10][234] = 35'b00000011111011111110011001011000000;
filter5[10][235] = 35'b00000001000000101100001011111100000;
filter5[10][236] = 35'b11111111000011100101101111101100000;
filter5[10][237] = 35'b00000000011001000010100110101001000;
filter5[10][238] = 35'b11111110111010111110001010110010000;
filter5[10][239] = 35'b11111111010110100001111001000110000;
filter5[10][240] = 35'b11111100001010010011101101100000000;
filter5[10][241] = 35'b00000000110100100100111011100100000;
filter5[10][242] = 35'b00000000100101011001000101101001000;
filter5[10][243] = 35'b00000000100001001011110010110010000;
filter5[10][244] = 35'b11111011000100111010010101111000000;
filter5[10][245] = 35'b00000010101110101101110100111100000;
filter5[10][246] = 35'b11111111001011001000111110011010000;
filter5[10][247] = 35'b00000000111010110010110110101110000;
filter5[10][248] = 35'b00000001101101000100111001011000000;
filter5[10][249] = 35'b00000100100110101101100000100000000;
filter5[10][250] = 35'b11111111111111101010101111000001000;
filter5[10][251] = 35'b00000010110101110100010110011100000;
filter5[10][252] = 35'b11111101101010010111011100001000000;
filter5[10][253] = 35'b00000001100001010011010111000100000;
filter5[10][254] = 35'b00000010101100100100100001010000000;
filter5[10][255] = 35'b00000001011101001011000001101000000;
filter5[10][256] = 35'b00000010000110111011100101110000000;
filter5[10][257] = 35'b00001000100000100111111111100000000;
filter5[10][258] = 35'b00001001000110011100011111110000000;
filter5[10][259] = 35'b11111011001111000001111011100000000;
filter5[10][260] = 35'b11110101100010101111001010010000000;
filter5[10][261] = 35'b11110111001110010000111001100000000;
filter5[10][262] = 35'b11110100011011011001010101110000000;
filter5[10][263] = 35'b11111101010010010100111000101000000;
filter5[10][264] = 35'b00001110000000111011000100100000000;
filter5[10][265] = 35'b00001011110001100010110001000000000;
filter5[10][266] = 35'b00000010100101101010010101110000000;
filter5[10][267] = 35'b11111000001110110100111101110000000;
filter5[10][268] = 35'b11111101110111001001110001100100000;
filter5[10][269] = 35'b00000100111000001100111001111000000;
filter5[10][270] = 35'b11111111101011100011101110110110100;
filter5[10][271] = 35'b11111011011110100011011101101000000;
filter5[10][272] = 35'b11111111000011111110100001100001000;
filter5[10][273] = 35'b11110110000010101110101010010000000;
filter5[10][274] = 35'b00000001111011111101111010000010000;
filter5[10][275] = 35'b11111111001011000001111010001010000;
filter5[10][276] = 35'b00000010011001010001000001000100000;
filter5[10][277] = 35'b00000001000001011010010110101100000;
filter5[10][278] = 35'b11111010011111110101110001011000000;
filter5[10][279] = 35'b11111001011111011011111000000000000;
filter5[10][280] = 35'b11111111101001000111100011101011000;
filter5[10][281] = 35'b11111001011000010000100000010000000;
filter5[10][282] = 35'b11111101100110011100111111001100000;
filter5[10][283] = 35'b11111101100110010100110110000000000;
filter5[10][284] = 35'b11111011001111100011110100110000000;
filter5[10][285] = 35'b11111100100011001000011001100000000;
filter5[10][286] = 35'b11111111000110100101001000010001000;
filter5[10][287] = 35'b00000011011100010101100110001100000;
filter5[10][288] = 35'b00000101011110001101100101111000000;
filter5[10][289] = 35'b11111100100111011000111101100000000;
filter5[10][290] = 35'b00000101010001101100011110001000000;
filter5[10][291] = 35'b00000000011110010110010101011010100;
filter5[10][292] = 35'b00000000011101011000011110101101100;
filter5[10][293] = 35'b11111110001000111110010010110100000;
filter5[10][294] = 35'b00000101111001100010011111101000000;
filter5[10][295] = 35'b00000011111101011101000010111100000;
filter5[10][296] = 35'b00000000101110110001001110000001000;
filter5[10][297] = 35'b11111111001001010001111001101111000;
filter5[10][298] = 35'b00000001100001101010011110111100000;
filter5[10][299] = 35'b11111111101011001001000101000111100;
filter5[10][300] = 35'b11111110101001101100001110011100000;
filter5[10][301] = 35'b00000010100000111000001000011000000;
filter5[10][302] = 35'b11111110101110101100100000100110000;
filter5[10][303] = 35'b00000011011111100101101010111000000;
filter5[10][304] = 35'b00000010100010010111110100111000000;
filter5[10][305] = 35'b11110111010000011001001010110000000;
filter5[10][306] = 35'b11111111001100011010111000100111000;
filter5[10][307] = 35'b11111111000010010000110010010001000;
filter5[10][308] = 35'b11111011101011000010100001110000000;
filter5[10][309] = 35'b11111111111101010011111100011101000;
filter5[10][310] = 35'b11111001011000011100100010110000000;
filter5[10][311] = 35'b00000001111000100101000000010100000;
filter5[10][312] = 35'b11111100101110001110010011100000000;
filter5[10][313] = 35'b11111100001010111010110110100100000;
filter5[10][314] = 35'b00000010100111000111011111100100000;
filter5[10][315] = 35'b00000010110110110110110000010100000;
filter5[10][316] = 35'b11111111000110001000001011011111000;
filter5[10][317] = 35'b00001000110111000010001111110000000;
filter5[10][318] = 35'b00000011001111010010001000101100000;
filter5[10][319] = 35'b11111011000100101000010111001000000;
filter5[10][320] = 35'b11111111101000001110100100000010100;
filter5[10][321] = 35'b00001011100010001011110110010000000;
filter5[10][322] = 35'b00000001001001001110111111111000000;
filter5[10][323] = 35'b11111010000101110101110111101000000;
filter5[10][324] = 35'b11110101101111000111010111110000000;
filter5[10][325] = 35'b11111100110011110010011111100100000;
filter5[10][326] = 35'b11111110111010010000001010101100000;
filter5[10][327] = 35'b11110010001111011000110000010000000;
filter5[10][328] = 35'b00000111100101000000100010011000000;
filter5[10][329] = 35'b11111110100001010001111100010110000;
filter5[10][330] = 35'b11111110011000110111100011100000000;
filter5[10][331] = 35'b11111000000110111111111001110000000;
filter5[10][332] = 35'b11111111011010111000000000101011000;
filter5[10][333] = 35'b00000001101011101111001011110110000;
filter5[10][334] = 35'b11111100111101110111000010110000000;
filter5[10][335] = 35'b11111110011111100011011011101010000;
filter5[10][336] = 35'b11111111111111011111000111010111001;
filter5[10][337] = 35'b00000000100011101100000101010000000;
filter5[10][338] = 35'b11111111111011111001001011001111101;
filter5[10][339] = 35'b11111111111000101001110110011001011;
filter5[10][340] = 35'b00000000111000111101110100101001000;
filter5[10][341] = 35'b00000011110010110110110001010100000;
filter5[10][342] = 35'b11111101100100000011111111000000000;
filter5[10][343] = 35'b11111010111110010100011110001000000;
filter5[10][344] = 35'b00000000000001101100000111000001000;
filter5[10][345] = 35'b11111110111100111001100111001110000;
filter5[10][346] = 35'b00000000110000011011011000110011000;
filter5[10][347] = 35'b11111110000110000010011010010000000;
filter5[10][348] = 35'b11111110011110111000100010101010000;
filter5[10][349] = 35'b11111111101110001100000000000110100;
filter5[10][350] = 35'b11111111111001011000001000001011100;
filter5[10][351] = 35'b00000010010101011111000001101100000;
filter5[10][352] = 35'b00000000001100001011101010100011000;
filter5[10][353] = 35'b00000001000100011100110011111100000;
filter5[10][354] = 35'b00000000110000000100000100010100000;
filter5[10][355] = 35'b00000010000101111000101010100000000;
filter5[10][356] = 35'b11111110000111010000011001010100000;
filter5[10][357] = 35'b11111110110000111010001011001010000;
filter5[10][358] = 35'b00000011110001000111101010010100000;
filter5[10][359] = 35'b11111110011011110101101010110000000;
filter5[10][360] = 35'b00000001011101101010101100100010000;
filter5[10][361] = 35'b00000000010010010000110101000110000;
filter5[10][362] = 35'b11111110100011101100010001110110000;
filter5[10][363] = 35'b00000000000101100010101101101110101;
filter5[10][364] = 35'b00000000001100000110100110111100010;
filter5[10][365] = 35'b00000000010101110110101101101100100;
filter5[10][366] = 35'b11111101101001011010111110011100000;
filter5[10][367] = 35'b11111111101010110100011100101110000;
filter5[10][368] = 35'b00000000110000000101101100001110000;
filter5[10][369] = 35'b00000001110011000010101100010010000;
filter5[10][370] = 35'b11111010010010111000011111000000000;
filter5[10][371] = 35'b00000001011100011011000111001000000;
filter5[10][372] = 35'b11111101100011000110001111010100000;
filter5[10][373] = 35'b00000001110111010110001001100000000;
filter5[10][374] = 35'b11111110110101011110100101111100000;
filter5[10][375] = 35'b11111110101001110001111000000100000;
filter5[10][376] = 35'b00000011010111111000001101001000000;
filter5[10][377] = 35'b00000101000011111001111100111000000;
filter5[10][378] = 35'b11111010011011110110010111011000000;
filter5[10][379] = 35'b00000011100100101100101010000100000;
filter5[10][380] = 35'b00000001000111011011001101111100000;
filter5[10][381] = 35'b11111110001010011100100111000100000;
filter5[10][382] = 35'b00000101101100101011010111000000000;
filter5[10][383] = 35'b00000100111111000000111100010000000;
filter5[10][384] = 35'b11111110101010111011100001011000000;
filter5[10][385] = 35'b11111101011010111011110111100100000;
filter5[10][386] = 35'b11111100111010001110110101001100000;
filter5[10][387] = 35'b11111110100011110101011010110000000;
filter5[10][388] = 35'b00000001010001011110100100100000000;
filter5[10][389] = 35'b11111101010010001010010111111100000;
filter5[10][390] = 35'b00000000000001111111010101001010101;
filter5[10][391] = 35'b00000010100001110101001110001000000;
filter5[10][392] = 35'b00000000010101010111101011100111100;
filter5[10][393] = 35'b11111100100111100001110110101100000;
filter5[10][394] = 35'b11111101001010100000111011101100000;
filter5[10][395] = 35'b00000000110000000111000000010010000;
filter5[10][396] = 35'b00000001001111111101000011100010000;
filter5[10][397] = 35'b00000100001000010110011011101000000;
filter5[10][398] = 35'b11111111110000111011111101100010100;
filter5[10][399] = 35'b11111111111100111010101101110010100;
filter5[10][400] = 35'b11111111111011010100011111010111111;
filter5[10][401] = 35'b11111111011011001000011011011011000;
filter5[10][402] = 35'b00000010010001000011000111001100000;
filter5[10][403] = 35'b00000000001011001001000101001110000;
filter5[10][404] = 35'b00000011011101111101011111101000000;
filter5[10][405] = 35'b00000000010100111100000010010010000;
filter5[10][406] = 35'b00000010100110100010011101000100000;
filter5[10][407] = 35'b11111100110000010111110011000100000;
filter5[10][408] = 35'b11111101001011101000111001100000000;
filter5[10][409] = 35'b00000001010011110110111100111010000;
filter5[10][410] = 35'b00000011100100010001101010011100000;
filter5[10][411] = 35'b00000100011111010011101100010000000;
filter5[10][412] = 35'b11111001101010100110001110111000000;
filter5[10][413] = 35'b00000011100000011110101110111000000;
filter5[10][414] = 35'b00000000001101100110010010110110110;
filter5[10][415] = 35'b11111110101001000000101000001100000;
filter5[10][416] = 35'b11111010010000001111110001011000000;
filter5[10][417] = 35'b00000000010001101010011101011000000;
filter5[10][418] = 35'b00000000100011010011011001010110000;
filter5[10][419] = 35'b00000000101001110101100000100010000;
filter5[10][420] = 35'b11111110000011110110110010010010000;
filter5[10][421] = 35'b11111101111000000010111010001000000;
filter5[10][422] = 35'b11111100111110101010111011001000000;
filter5[10][423] = 35'b11111111111110010100001010001011011;
filter5[10][424] = 35'b11111110011001101111111110000110000;
filter5[10][425] = 35'b11111110100110001011100011111100000;
filter5[10][426] = 35'b00000000001111001101110001001111110;
filter5[10][427] = 35'b11111101010001100110100101100100000;
filter5[10][428] = 35'b00000000110100010100000100100101000;
filter5[10][429] = 35'b11111110001101111110010101010000000;
filter5[10][430] = 35'b00000000000000100000001100101000111;
filter5[10][431] = 35'b00000000010110111101100000010001100;
filter5[10][432] = 35'b11110100100100000000000000010000000;
filter5[10][433] = 35'b00000011010110100100000100110000000;
filter5[10][434] = 35'b00000000101000011011111000100001000;
filter5[10][435] = 35'b11111011110110110010001111011000000;
filter5[10][436] = 35'b00000000011010111011111100000110000;
filter5[10][437] = 35'b00000000100011100011010110001000000;
filter5[10][438] = 35'b00000001111011101100100011001110000;
filter5[10][439] = 35'b00000000111110101011010011000100000;
filter5[10][440] = 35'b00000001011100011110010001010100000;
filter5[10][441] = 35'b11111001101110001010100010011000000;
filter5[10][442] = 35'b00000011010000101111100111011000000;
filter5[10][443] = 35'b11111000111110011001110011111000000;
filter5[10][444] = 35'b00000101011000110111111010010000000;
filter5[10][445] = 35'b00000000100111011010000000110110000;
filter5[10][446] = 35'b11111101010001010010100100111000000;
filter5[10][447] = 35'b11111111010111000001011111000001000;
filter5[10][448] = 35'b11111101010001011011100011101000000;
filter5[10][449] = 35'b11110100001000010010001000010000000;
filter5[10][450] = 35'b11110011000011000011101101110000000;
filter5[10][451] = 35'b11111000001100100011100111001000000;
filter5[10][452] = 35'b11111110100001111001111101000010000;
filter5[10][453] = 35'b11111011010011111010000001000000000;
filter5[10][454] = 35'b00000000101011110001111001001101000;
filter5[10][455] = 35'b00000000011101101110101000100010100;
filter5[10][456] = 35'b11111000111100011101111001000000000;
filter5[10][457] = 35'b00000000001000110011110110110101100;
filter5[10][458] = 35'b00000010111100101011011001011000000;
filter5[10][459] = 35'b00000100010011110111010000000000000;
filter5[10][460] = 35'b00000111010111100000100100011000000;
filter5[10][461] = 35'b00000111000111100010110111100000000;
filter5[10][462] = 35'b00000000101101010110101001111011000;
filter5[10][463] = 35'b00000011101100011011000001111100000;
filter5[10][464] = 35'b11111011100011010010011100100000000;
filter5[10][465] = 35'b00000100001101010011100011101000000;
filter5[10][466] = 35'b00010010111111111110101101000000000;
filter5[10][467] = 35'b00010000101101010100100110000000000;
filter5[10][468] = 35'b00010101100010111011000000000000000;
filter5[10][469] = 35'b00000011110011100111001100000000000;
filter5[10][470] = 35'b11111111011101011110000001011110000;
filter5[10][471] = 35'b11111001110100111100011110001000000;
filter5[10][472] = 35'b00000000100000101000100111110001000;
filter5[10][473] = 35'b11111110001100001001010000011000000;
filter5[10][474] = 35'b00001010010101100101000001010000000;
filter5[10][475] = 35'b11111111110100001100111111111111100;
filter5[10][476] = 35'b11111100111100101111011010111100000;
filter5[10][477] = 35'b11111110011000101011011111011010000;
filter5[10][478] = 35'b00000010001011011100010111101000000;
filter5[10][479] = 35'b11110111001000111111001010110000000;
filter5[10][480] = 35'b11111001011111010011100101110000000;
filter5[10][481] = 35'b11111011001101101100101001100000000;
filter5[10][482] = 35'b00000010001100000011100011010100000;
filter5[10][483] = 35'b11111011111011110110110111100000000;
filter5[10][484] = 35'b11111011101110001010001101101000000;
filter5[10][485] = 35'b11111110011010000111010010010000000;
filter5[10][486] = 35'b11111101111001010110011101001100000;
filter5[10][487] = 35'b11111010110101101001011111010000000;
filter5[10][488] = 35'b00000010110111101001101000000000000;
filter5[10][489] = 35'b00000010011011110000001110000100000;
filter5[10][490] = 35'b00001000101000100000000100110000000;
filter5[10][491] = 35'b11110100111100011111101111100000000;
filter5[10][492] = 35'b11111011111010111010111010000000000;
filter5[10][493] = 35'b00000110110100001001101110100000000;
filter5[10][494] = 35'b00000001100010000111110100010000000;
filter5[10][495] = 35'b00000001110010000000100001101000000;
filter5[10][496] = 35'b00000010001101010000111111010000000;
filter5[10][497] = 35'b00000011110100011100100110011100000;
filter5[10][498] = 35'b11111111110010101110001101110011000;
filter5[10][499] = 35'b11111101100110001100001110001100000;
filter5[10][500] = 35'b11111110110100001111100001101010000;
filter5[10][501] = 35'b00000000001001000001000100000111100;
filter5[10][502] = 35'b00000010100101110101100010100000000;
filter5[10][503] = 35'b00000000001101101100011110111110010;
filter5[10][504] = 35'b00000011011100110111000010111100000;
filter5[10][505] = 35'b11111110111100101010101011011000000;
filter5[10][506] = 35'b00000110100111101011001011110000000;
filter5[10][507] = 35'b11111010101011110110010101111000000;
filter5[10][508] = 35'b11111010010011101100110101111000000;
filter5[10][509] = 35'b00000000110001100110111001100001000;
filter5[10][510] = 35'b00000100010011001101101010010000000;
filter5[10][511] = 35'b11111101100111110010010101000100000;
filter5[10][512] = 35'b11111001011110110101110110110000000;
filter5[10][513] = 35'b00000011001100001010101001010000000;
filter5[10][514] = 35'b00000001001000111011101001001010000;
filter5[10][515] = 35'b00000010010101011000011100101100000;
filter5[10][516] = 35'b11111100101011100010001101010100000;
filter5[10][517] = 35'b00000001111011010011110111101100000;
filter5[10][518] = 35'b11111110000010100100000011001110000;
filter5[10][519] = 35'b11111011000001110110100010110000000;
filter5[10][520] = 35'b00000000110111011011010101001101000;
filter5[10][521] = 35'b11111110100010110000010101110000000;
filter5[10][522] = 35'b00000000111101011001010011101010000;
filter5[10][523] = 35'b00000011011011001110000110100000000;
filter5[10][524] = 35'b11111110000100001001101100001110000;
filter5[10][525] = 35'b11111111011100100011100100010111000;
filter5[10][526] = 35'b11111110110101011010000011000010000;
filter5[10][527] = 35'b11111101010101111001010010101000000;
filter5[10][528] = 35'b00000011101001001000011011100100000;
filter5[10][529] = 35'b00000001001010010100101111110010000;
filter5[10][530] = 35'b11111110111110011101111011010110000;
filter5[10][531] = 35'b00000000111010110101111100000100000;
filter5[10][532] = 35'b00000011100101001110110101111000000;
filter5[10][533] = 35'b11111111010100011010000111001011000;
filter5[10][534] = 35'b11111111010010100001101001101110000;
filter5[10][535] = 35'b11111110001001110101101010001100000;
filter5[10][536] = 35'b00000000101001010110001100100101000;
filter5[10][537] = 35'b00000001011110101011100110111010000;
filter5[10][538] = 35'b11111101111110101101001111010000000;
filter5[10][539] = 35'b00000010000001111111010010001000000;
filter5[10][540] = 35'b11111101001010000000100001110100000;
filter5[10][541] = 35'b00000011110011010010000101000000000;
filter5[10][542] = 35'b00000001110101001001100110101110000;
filter5[10][543] = 35'b11111111010100110000010100101110000;
filter5[10][544] = 35'b11111011010000010011010000101000000;
filter5[10][545] = 35'b11111111110101001101011001110111010;
filter5[10][546] = 35'b00000010101010111111011010001000000;
filter5[10][547] = 35'b11111011011010111011100001000000000;
filter5[10][548] = 35'b11111111001101111011100000011001000;
filter5[10][549] = 35'b00000100011011010011110001100000000;
filter5[10][550] = 35'b11111111001100001001110001001010000;
filter5[10][551] = 35'b11111111000001111010101101111101000;
filter5[10][552] = 35'b00000010010110011000000000011000000;
filter5[10][553] = 35'b11111111010110110000110011001100000;
filter5[10][554] = 35'b00000010100011100101111010011100000;
filter5[10][555] = 35'b11111111000111001011101110110100000;
filter5[10][556] = 35'b00000000001001000100100010101111100;
filter5[10][557] = 35'b11111100110000101001000011101000000;
filter5[10][558] = 35'b00000011010010100000100001100000000;
filter5[10][559] = 35'b11111111011111110110100010001100000;
filter5[10][560] = 35'b11111101110011101111111001110000000;
filter5[10][561] = 35'b11111111010100000111100010100111000;
filter5[10][562] = 35'b11111101001000000010101110101000000;
filter5[10][563] = 35'b00000010101110011101100011010000000;
filter5[10][564] = 35'b11111111001100001000011100001101000;
filter5[10][565] = 35'b11111011110110111100100101001000000;
filter5[10][566] = 35'b11111110111111100000000111000010000;
filter5[10][567] = 35'b11111100010101011111000100101100000;
filter5[10][568] = 35'b00000001100110010111011111011000000;
filter5[10][569] = 35'b00000011010100010011110011001000000;
filter5[10][570] = 35'b00000000110100101100100000010011000;
filter5[10][571] = 35'b11111111111111110101000101010001100;
filter5[10][572] = 35'b00000001011101100011000110011000000;
filter5[10][573] = 35'b11111111000010010100111010111100000;
filter5[10][574] = 35'b11111110111010110000011010101010000;
filter5[10][575] = 35'b00000011000011011001101010101000000;
filter5[10][576] = 35'b11111011111101101101110100100000000;
filter5[10][577] = 35'b00000010000101111100011110100100000;
filter5[10][578] = 35'b00000010010110110001010110011100000;
filter5[10][579] = 35'b00000000111001111010010101010100000;
filter5[10][580] = 35'b11111010010101100101101000011000000;
filter5[10][581] = 35'b11111111111011110010001000100101111;
filter5[10][582] = 35'b11111100001011110010100001010000000;
filter5[10][583] = 35'b11111010110110100010111010011000000;
filter5[10][584] = 35'b11110111110000011100000011100000000;
filter5[10][585] = 35'b00000101110011011110010100000000000;
filter5[10][586] = 35'b00000010100011010000101010010000000;
filter5[10][587] = 35'b00000010001001111110011011100000000;
filter5[10][588] = 35'b11111111000110100110111111010111000;
filter5[10][589] = 35'b00000011011001001101001111001000000;
filter5[10][590] = 35'b11111101101101001001010010010000000;
filter5[10][591] = 35'b11111111111110001100110000001010001;
filter5[10][592] = 35'b11111111011001101110011001111011000;
filter5[10][593] = 35'b00000010010100011010110001111000000;
filter5[10][594] = 35'b00000011100000000010010110111100000;
filter5[10][595] = 35'b00000000001010100010001010110111010;
filter5[10][596] = 35'b00000010010010111000100100000000000;
filter5[10][597] = 35'b00000001010100010000011111001100000;
filter5[10][598] = 35'b11111111110011011000110010100111010;
filter5[10][599] = 35'b11111110101010111001000000000000000;
filter5[10][600] = 35'b11111100001001010110101011000000000;
filter5[10][601] = 35'b11111100010011010000000100100000000;
filter5[10][602] = 35'b00000010101010111111000110100100000;
filter5[10][603] = 35'b11111010001001010011101000000000000;
filter5[10][604] = 35'b11111101000001011111101101101000000;
filter5[10][605] = 35'b00000000001101010001100001101100100;
filter5[10][606] = 35'b00000100000100001110010111110000000;
filter5[10][607] = 35'b11111010100011011001110110000000000;
filter5[10][608] = 35'b11111001000001001101000000011000000;
filter5[10][609] = 35'b00000000000100100000100000000101111;
filter5[10][610] = 35'b11111101111010000001010100010000000;
filter5[10][611] = 35'b00000010101101000001000011011000000;
filter5[10][612] = 35'b11111100011101100101010101111000000;
filter5[10][613] = 35'b00000000010000101110011010001000000;
filter5[10][614] = 35'b11111111111001000111011010010111110;
filter5[10][615] = 35'b11111111111011000101100010000000101;
filter5[10][616] = 35'b11111111000000111100011000101010000;
filter5[10][617] = 35'b00000000000100111011001101111100111;
filter5[10][618] = 35'b11111100101001111011010001111000000;
filter5[10][619] = 35'b00000011001011100010110001000100000;
filter5[10][620] = 35'b00000000000010001010110011111010100;
filter5[10][621] = 35'b11111111011010001100110101101110000;
filter5[10][622] = 35'b11111111010101111100001110101011000;
filter5[10][623] = 35'b11111101000010111111001110010000000;
filter5[10][624] = 35'b00000000101011001010100101111010000;
filter5[10][625] = 35'b00000000001111000011011001111111010;
filter5[10][626] = 35'b11111101101010010010001001010100000;
filter5[10][627] = 35'b11111111010000111110101000110000000;
filter5[10][628] = 35'b11111101100110001000001011011000000;
filter5[10][629] = 35'b11111111011111111000000010100001000;
filter5[10][630] = 35'b11111111011000110110010000010111000;
filter5[10][631] = 35'b00000000011101100101100111101000000;
filter5[10][632] = 35'b00000101000110100001011111001000000;
filter5[10][633] = 35'b11111110000111011111101110010100000;
filter5[10][634] = 35'b00000010101101101100101100110000000;
filter5[10][635] = 35'b11111111100001000100101010011011000;
filter5[10][636] = 35'b11111111101001000100111110011110100;
filter5[10][637] = 35'b00000000100001001110011100011110000;
filter5[10][638] = 35'b00000101001111001101111001100000000;
filter5[10][639] = 35'b00000001011111101000101000101100000;
filter5[10][640] = 35'b11110011101111110011101011100000000;
filter5[10][641] = 35'b11111011110100010001101001001000000;
filter5[10][642] = 35'b11111110111000001111000111100010000;
filter5[10][643] = 35'b00000101100000000000011011111000000;
filter5[10][644] = 35'b11111111110001110100101100110000100;
filter5[10][645] = 35'b00000010010000011101001101111100000;
filter5[10][646] = 35'b00000110101101100100110011001000000;
filter5[10][647] = 35'b00000011111111101000001100110000000;
filter5[10][648] = 35'b11111001001111111000010010110000000;
filter5[10][649] = 35'b11111011011000110100110100001000000;
filter5[10][650] = 35'b00000011111011001110101111000000000;
filter5[10][651] = 35'b00000101010011100001101000100000000;
filter5[10][652] = 35'b00000000110011100111100010001010000;
filter5[10][653] = 35'b11111110010110001101110110011010000;
filter5[10][654] = 35'b00000000100110011111010001001000000;
filter5[10][655] = 35'b00000000101000010110110011000011000;
filter5[10][656] = 35'b11111100101000110100010100100100000;
filter5[10][657] = 35'b00001100110111011010011110010000000;
filter5[10][658] = 35'b00001111001010000001010000010000000;
filter5[10][659] = 35'b00001010010011101100001111100000000;
filter5[10][660] = 35'b00000001110100110010101101001100000;
filter5[10][661] = 35'b00000000100110001111101001101110000;
filter5[10][662] = 35'b11111110110111011000010010010000000;
filter5[10][663] = 35'b11111000100111001011000100010000000;
filter5[10][664] = 35'b11111111011010101000011001011000000;
filter5[10][665] = 35'b11111101101001010011100000111100000;
filter5[10][666] = 35'b00000110111010100001000000011000000;
filter5[10][667] = 35'b11111100100110000011000000111000000;
filter5[10][668] = 35'b00000100000101010100010011011000000;
filter5[10][669] = 35'b11111110010010110000100010110000000;
filter5[10][670] = 35'b11111110011011110111000101011010000;
filter5[10][671] = 35'b11111110111011100100101000111110000;
filter5[10][672] = 35'b11111001100011101101110000011000000;
filter5[10][673] = 35'b11111010000000110110110011111000000;
filter5[10][674] = 35'b11111111100100000110001010111010000;
filter5[10][675] = 35'b00000000110110000101100010011111000;
filter5[10][676] = 35'b11111001110111101001010110110000000;
filter5[10][677] = 35'b11111101001000010100001000001000000;
filter5[10][678] = 35'b00000000000000111010100110000110100;
filter5[10][679] = 35'b11111100001010110000010011111100000;
filter5[10][680] = 35'b00000011101100011000011011001000000;
filter5[10][681] = 35'b00000011111000001000100011010100000;
filter5[10][682] = 35'b11111111100010011111010110000010100;
filter5[10][683] = 35'b11111100100100101010111111001000000;
filter5[10][684] = 35'b11111111000111101110101010110001000;
filter5[10][685] = 35'b11111111011100110110011100001111000;
filter5[10][686] = 35'b00000000011101010101111101000000000;
filter5[10][687] = 35'b00000011011100000001101110111000000;
filter5[10][688] = 35'b00000001010000000101111110100000000;
filter5[10][689] = 35'b11111110011100110011110001111110000;
filter5[10][690] = 35'b11111101000100101001001110111000000;
filter5[10][691] = 35'b11111110100010001010001001101010000;
filter5[10][692] = 35'b00000010010110100011000101000000000;
filter5[10][693] = 35'b00000000110001101100001111010110000;
filter5[10][694] = 35'b00000001000001110001111000110110000;
filter5[10][695] = 35'b11111101001001101111101000110000000;
filter5[10][696] = 35'b11111101100011000111000001101100000;
filter5[10][697] = 35'b00000010110101011110110011000100000;
filter5[10][698] = 35'b00000001011101101001000110000000000;
filter5[10][699] = 35'b11111100010111110100001011101000000;
filter5[10][700] = 35'b00000010010110111101101010011000000;
filter5[10][701] = 35'b00000001010110010101111110100000000;
filter5[10][702] = 35'b00000000011100110111100010011010100;
filter5[10][703] = 35'b00000000100011101101101100011100000;
filter5[10][704] = 35'b11111111111100001111001111011001110;
filter5[10][705] = 35'b00000010010111100011100110100100000;
filter5[10][706] = 35'b11111111011011000011101000111100000;
filter5[10][707] = 35'b00000000100011110011111101000111000;
filter5[10][708] = 35'b11111111010000111000010011010011000;
filter5[10][709] = 35'b00000000101001110001111100011011000;
filter5[10][710] = 35'b00000000001100011101101001000100110;
filter5[10][711] = 35'b11111111001001011111011110011101000;
filter5[10][712] = 35'b00000010101001110101001101101000000;
filter5[10][713] = 35'b00000000100110011111101111001000000;
filter5[10][714] = 35'b11111111011101101011101111101110000;
filter5[10][715] = 35'b11111111000111010111100010011101000;
filter5[10][716] = 35'b00000001101000101001000011101010000;
filter5[10][717] = 35'b00000001000101101111010100111110000;
filter5[10][718] = 35'b11111111110101111101110110100000000;
filter5[10][719] = 35'b11111110111010000010100100000000000;
filter5[10][720] = 35'b00000001111101000010111000010110000;
filter5[10][721] = 35'b11111111100111001101001001111011100;
filter5[10][722] = 35'b11111110010101000100001110010100000;
filter5[10][723] = 35'b00000010000010010100000100010100000;
filter5[10][724] = 35'b00000001001001101111110000001000000;
filter5[10][725] = 35'b00000010000111010000101110010100000;
filter5[10][726] = 35'b11111100010111100110110000101100000;
filter5[10][727] = 35'b11111111110111001101101100111011100;
filter5[10][728] = 35'b11111111000100001000100100000001000;
filter5[10][729] = 35'b11111011001100110000010101010000000;
filter5[10][730] = 35'b00000000000011001100101111010011010;
filter5[10][731] = 35'b00000000100111011000101110011111000;
filter5[10][732] = 35'b00000000110000100011101100000000000;
filter5[10][733] = 35'b00000000010101100111111100100111000;
filter5[10][734] = 35'b11111110000010100011010111110010000;
filter5[10][735] = 35'b00000000010110100101011100000001000;
filter5[10][736] = 35'b00000001110010011101110000110100000;
filter5[10][737] = 35'b11111100100010101100011110101000000;
filter5[10][738] = 35'b00000011011011000000011101111100000;
filter5[10][739] = 35'b11111100111001110010101000001100000;
filter5[10][740] = 35'b11111101101110101111110111110100000;
filter5[10][741] = 35'b11111101010111101100110110100100000;
filter5[10][742] = 35'b00000100110001110011000110111000000;
filter5[10][743] = 35'b00000000010110111111101001100101100;
filter5[10][744] = 35'b11111111001101001000100011101100000;
filter5[10][745] = 35'b00000010010000101110011110110000000;
filter5[10][746] = 35'b00000001100110101011111100110010000;
filter5[10][747] = 35'b11111101011101110000101111111100000;
filter5[10][748] = 35'b11111101011000001010000011110100000;
filter5[10][749] = 35'b00000001110110100000010000111100000;
filter5[10][750] = 35'b11111110000110010100010111000010000;
filter5[10][751] = 35'b11111111001000001110110011101110000;
filter5[10][752] = 35'b00000000000001010110100000100001101;
filter5[10][753] = 35'b00000011110101010110111011101100000;
filter5[10][754] = 35'b11111101011110111010001010110000000;
filter5[10][755] = 35'b00000000010000000011001011111110100;
filter5[10][756] = 35'b11111111001111110010111111110010000;
filter5[10][757] = 35'b00000010110011001101010100100000000;
filter5[10][758] = 35'b11111110001001000101100101010100000;
filter5[10][759] = 35'b00000010101011001111101000010100000;
filter5[10][760] = 35'b00000000101100101100011010000111000;
filter5[10][761] = 35'b00000101110001100010011001010000000;
filter5[10][762] = 35'b00000010011001010001001010110000000;
filter5[10][763] = 35'b00000001001111011010111011110010000;
filter5[10][764] = 35'b11111101010110011010000101110000000;
filter5[10][765] = 35'b00000011111100011101111000101000000;
filter5[10][766] = 35'b00000000100111000110011101110010000;
filter5[10][767] = 35'b11111100110011011011010111110100000;
filter5[10][768] = 35'b11111111000011110010111010101000000;
filter5[10][769] = 35'b11111001110001101101011000000000000;
filter5[10][770] = 35'b11111000100110011000001101011000000;
filter5[10][771] = 35'b00000000101000111011111111111110000;
filter5[10][772] = 35'b11111111100101100000111100110110000;
filter5[10][773] = 35'b00000010010100000100010001001100000;
filter5[10][774] = 35'b00000001000010000001100000110110000;
filter5[10][775] = 35'b11111101011000110011000010101100000;
filter5[10][776] = 35'b11111001001101101100100101000000000;
filter5[10][777] = 35'b11110110111111011101100100010000000;
filter5[10][778] = 35'b00001001010111011001011000000000000;
filter5[10][779] = 35'b11111110010011001100101010110010000;
filter5[10][780] = 35'b00000100000000100101111100100000000;
filter5[10][781] = 35'b11111110000110011010001001101110000;
filter5[10][782] = 35'b11111111100000010100111000011110000;
filter5[10][783] = 35'b11111111111010010001011001101101000;
filter5[10][784] = 35'b11111011110001001101010100010000000;
filter5[10][785] = 35'b11111101010111111101100001110100000;
filter5[10][786] = 35'b00001010010000011101001111010000000;
filter5[10][787] = 35'b00000001111100111010000011101110000;
filter5[10][788] = 35'b00000110010100111010000100011000000;
filter5[10][789] = 35'b00000011110101010011001010100000000;
filter5[10][790] = 35'b00000100101011000100010011001000000;
filter5[10][791] = 35'b00000010010110111000001100010000000;
filter5[10][792] = 35'b11111111100111011001101100011011000;
filter5[10][793] = 35'b00000000001010111001100011111111100;
filter5[10][794] = 35'b00000001101011011010000100001110000;
filter5[10][795] = 35'b00000110010100000101000111010000000;
filter5[10][796] = 35'b11111110010010000010011001000110000;
filter5[10][797] = 35'b00000011011011000010001100011100000;
filter5[10][798] = 35'b00000101000111101000011000111000000;
filter5[10][799] = 35'b11111111110110100110110011101111110;
filter5[10][800] = 35'b11111101111011101111010011000000000;
filter5[10][801] = 35'b00000001011111010010011101011110000;
filter5[10][802] = 35'b11111101011010111000110010110000000;
filter5[10][803] = 35'b11111111011110111111001110110110000;
filter5[10][804] = 35'b11111101001000111010001010100000000;
filter5[10][805] = 35'b11111101110001101000000000111100000;
filter5[10][806] = 35'b11111100010011100100010100000000000;
filter5[10][807] = 35'b11111010110101011100001001101000000;
filter5[10][808] = 35'b11111101100110111110001100001000000;
filter5[10][809] = 35'b00000000011101010101010111001001000;
filter5[10][810] = 35'b11111101101010010010110011001100000;
filter5[10][811] = 35'b11111101000110101001001001000100000;
filter5[10][812] = 35'b11111111000110100000110100000001000;
filter5[10][813] = 35'b00000000111011111110101101100010000;
filter5[10][814] = 35'b11111101110101101010111101111000000;
filter5[10][815] = 35'b11111111010101111011110111001010000;
filter5[10][816] = 35'b00000010000001110010000111100100000;
filter5[10][817] = 35'b00000101000101101000001100000000000;
filter5[10][818] = 35'b11111111001101101110110101001000000;
filter5[10][819] = 35'b00000011000100110101010111010000000;
filter5[10][820] = 35'b00000001101111100010110011001010000;
filter5[10][821] = 35'b00000000001010001001101010101100100;
filter5[10][822] = 35'b00000010101110111100111111001100000;
filter5[10][823] = 35'b11111110101111011100100110010100000;
filter5[10][824] = 35'b00000001010010000001011100110000000;
filter5[10][825] = 35'b11111111010111111111011011011100000;
filter5[10][826] = 35'b11111000100100101100010000000000000;
filter5[10][827] = 35'b00000100111001110110001111110000000;
filter5[10][828] = 35'b11111100100111000111001011010100000;
filter5[10][829] = 35'b11111100010101100101100101000000000;
filter5[10][830] = 35'b00000010110010110110101110010000000;
filter5[10][831] = 35'b11111111110010001111101101101011010;
filter5[10][832] = 35'b00000000101011111110111111000000000;
filter5[10][833] = 35'b00000000100101100001100101110100000;
filter5[10][834] = 35'b00000001010010110111011110110000000;
filter5[10][835] = 35'b00000000101010010100001010000101000;
filter5[10][836] = 35'b00000000001100011110000101110101000;
filter5[10][837] = 35'b11111111111101100100100110111010010;
filter5[10][838] = 35'b11111111100010000110001010101011000;
filter5[10][839] = 35'b11111111100000110011000100110010000;
filter5[10][840] = 35'b11111111011010100110001101000011000;
filter5[10][841] = 35'b00000001101000010110010001000110000;
filter5[10][842] = 35'b00000000000001001011000101110001010;
filter5[10][843] = 35'b00000001101111110000010100111010000;
filter5[10][844] = 35'b11111110011111101111110111000100000;
filter5[10][845] = 35'b00000000010000110010000001011001100;
filter5[10][846] = 35'b00000000110010110100011101001000000;
filter5[10][847] = 35'b11111111110001110101101010101000110;
filter5[10][848] = 35'b00000000110010101101111001100111000;
filter5[10][849] = 35'b11111111000110010000010001100000000;
filter5[10][850] = 35'b11111101100110010000001011011100000;
filter5[10][851] = 35'b00000011011101001011100111100100000;
filter5[10][852] = 35'b00000000111110111111111011110111000;
filter5[10][853] = 35'b00000010100010011011101111101000000;
filter5[10][854] = 35'b11111111010000010010001010010001000;
filter5[10][855] = 35'b11111111000000100001000110110000000;
filter5[10][856] = 35'b00000000101111101010100011010000000;
filter5[10][857] = 35'b11111111000000011001101101000001000;
filter5[10][858] = 35'b00000000001111011010100010111110110;
filter5[10][859] = 35'b11111100001010101100001010010000000;
filter5[10][860] = 35'b00000010101101001011001110110000000;
filter5[10][861] = 35'b00000001111011010110110011000110000;
filter5[10][862] = 35'b11111110111110010001100001001100000;
filter5[10][863] = 35'b00000000111001111111010101010101000;
filter5[10][864] = 35'b00000001010110100111011001011100000;
filter5[10][865] = 35'b11111100101100000010111111010100000;
filter5[10][866] = 35'b00000000000010101110101110110101100;
filter5[10][867] = 35'b00000000100011000011101000010011000;
filter5[10][868] = 35'b00000000100000111001111010010001000;
filter5[10][869] = 35'b11111110100110101100011111101110000;
filter5[10][870] = 35'b00000001101010111100000100001010000;
filter5[10][871] = 35'b00000011000111101110010000001100000;
filter5[10][872] = 35'b11111111101100101111110001011011100;
filter5[10][873] = 35'b11111110010111110010101110001100000;
filter5[10][874] = 35'b00000110100110001001011001100000000;
filter5[10][875] = 35'b11111111011111011010111010101010000;
filter5[10][876] = 35'b11111101001100111010110010101000000;
filter5[10][877] = 35'b11111110101110111101110100110010000;
filter5[10][878] = 35'b00000011001001000101001101100000000;
filter5[10][879] = 35'b00000010011010101100101110010100000;
filter5[10][880] = 35'b00000010101100111000010010000000000;
filter5[10][881] = 35'b11111100001010000001101101000000000;
filter5[10][882] = 35'b11111111001100001001011011110110000;
filter5[10][883] = 35'b11111100111111000011100110010100000;
filter5[10][884] = 35'b11111111011000000100001101101000000;
filter5[10][885] = 35'b00000001001000000110111110111010000;
filter5[10][886] = 35'b11111010000101010001001110000000000;
filter5[10][887] = 35'b00000000000010100110111111000101010;
filter5[10][888] = 35'b00000000001111100100110000111100010;
filter5[10][889] = 35'b11111111010000000101110101001011000;
filter5[10][890] = 35'b00000110000000001101101110100000000;
filter5[10][891] = 35'b11111100011111010010010101010100000;
filter5[10][892] = 35'b00000000011110111110001000101111000;
filter5[10][893] = 35'b00000101000101011010110001010000000;
filter5[10][894] = 35'b00000100110010111100000000010000000;
filter5[10][895] = 35'b00000000101011000011110101111110000;
filter5[10][896] = 35'b00000100101101011000101101111000000;
filter5[10][897] = 35'b00001000001010011110010001010000000;
filter5[10][898] = 35'b00000001000011101100011011011010000;
filter5[10][899] = 35'b11111010101010110101111001011000000;
filter5[10][900] = 35'b11111001010100010000110100011000000;
filter5[10][901] = 35'b11111101011100101001010111100000000;
filter5[10][902] = 35'b11111111010001101001100101001011000;
filter5[10][903] = 35'b11110100011111001100010101000000000;
filter5[10][904] = 35'b00001001100000100011110101000000000;
filter5[10][905] = 35'b11111101010110000110001110110000000;
filter5[10][906] = 35'b11111110000110010111011001000000000;
filter5[10][907] = 35'b00000001100101011001000001010110000;
filter5[10][908] = 35'b00000100011111110111010010011000000;
filter5[10][909] = 35'b00000010000101100111001100010000000;
filter5[10][910] = 35'b11111101100101010011110111011100000;
filter5[10][911] = 35'b11111100100111011010101100000000000;
filter5[10][912] = 35'b00000010011110001111110100000100000;
filter5[10][913] = 35'b00000000100001000101110011010111000;
filter5[10][914] = 35'b11111101100010010111000010011000000;
filter5[10][915] = 35'b00000100110011000111001001100000000;
filter5[10][916] = 35'b00000011000110011011011111000000000;
filter5[10][917] = 35'b00000001000000010010111000101100000;
filter5[10][918] = 35'b11111010010101101111001111011000000;
filter5[10][919] = 35'b11111111101011110111101100101110100;
filter5[10][920] = 35'b11111101100011101111101111101000000;
filter5[10][921] = 35'b11111010010100001110101011110000000;
filter5[10][922] = 35'b00000000010100001110011010100110000;
filter5[10][923] = 35'b11111100110011001001110100110000000;
filter5[10][924] = 35'b11111111001110101011011011110011000;
filter5[10][925] = 35'b00000001110111000100101000000010000;
filter5[10][926] = 35'b00000000000001011111011011000010010;
filter5[10][927] = 35'b00000101110001101101010111100000000;
filter5[10][928] = 35'b00000011010011010110011111010000000;
filter5[10][929] = 35'b11111010110111001011110111111000000;
filter5[10][930] = 35'b00000011001100001010011110110100000;
filter5[10][931] = 35'b11111111010000000110110110110011000;
filter5[10][932] = 35'b11111110101110000001100111111100000;
filter5[10][933] = 35'b11111100111010011001100001111100000;
filter5[10][934] = 35'b00000000101000111010110101001101000;
filter5[10][935] = 35'b00000100010110111001110001100000000;
filter5[10][936] = 35'b11111111011001011110110101011100000;
filter5[10][937] = 35'b00000001010000100000000010000000000;
filter5[10][938] = 35'b00000001000110001010111001111110000;
filter5[10][939] = 35'b00000000100011011101001010000100000;
filter5[10][940] = 35'b11111111001000110001101110111111000;
filter5[10][941] = 35'b00000001001101001000100010001000000;
filter5[10][942] = 35'b11111101110000111001110110111100000;
filter5[10][943] = 35'b00000010110111100010100010111000000;
filter5[10][944] = 35'b00000001101000101101111111011010000;
filter5[10][945] = 35'b00000001010111001100111000010000000;
filter5[10][946] = 35'b11111110101011100111001011100010000;
filter5[10][947] = 35'b11111100111000001110010111101100000;
filter5[10][948] = 35'b11111110101110011010111011101000000;
filter5[10][949] = 35'b00000101000001100100000101100000000;
filter5[10][950] = 35'b11111001100101010000010010111000000;
filter5[10][951] = 35'b00000011111001011111000011101100000;
filter5[10][952] = 35'b11111111111000011000100101001100111;
filter5[10][953] = 35'b00000011110001111100011011100000000;
filter5[10][954] = 35'b11111101110011100001100010101100000;
filter5[10][955] = 35'b00000001111001111110010110010100000;
filter5[10][956] = 35'b00000000101000000001100000101111000;
filter5[10][957] = 35'b00000001111001000000110101100100000;
filter5[10][958] = 35'b00001000111110111111110100110000000;
filter5[10][959] = 35'b00001011101100011001111000000000000;
filter5[10][960] = 35'b11111001101100101101010101100000000;
filter5[10][961] = 35'b00000101110010101011100111010000000;
filter5[10][962] = 35'b00000101000001000101101001010000000;
filter5[10][963] = 35'b00000001110000111110101101101110000;
filter5[10][964] = 35'b11111100000110000111011101110000000;
filter5[10][965] = 35'b11111011011000010110001110011000000;
filter5[10][966] = 35'b00000000001101001000011010001001110;
filter5[10][967] = 35'b11111100001101111101100101010000000;
filter5[10][968] = 35'b00000101110110101010010110111000000;
filter5[10][969] = 35'b11111111100100111000111100111011000;
filter5[10][970] = 35'b11111110101001101101100111001000000;
filter5[10][971] = 35'b11111111100110100100101110000000100;
filter5[10][972] = 35'b00000011100111111011101110101100000;
filter5[10][973] = 35'b00000010000100101001000100111100000;
filter5[10][974] = 35'b11111101110101000000100110001000000;
filter5[10][975] = 35'b00000000000111111010101101011101110;
filter5[10][976] = 35'b11111110111001010101000101001110000;
filter5[10][977] = 35'b11111110010010101100100110010010000;
filter5[10][978] = 35'b11111100111010010111010100011100000;
filter5[10][979] = 35'b11111111001010100010001001111010000;
filter5[10][980] = 35'b00000001101000011100100110110000000;
filter5[10][981] = 35'b00000010110011100010001010110100000;
filter5[10][982] = 35'b11111110101000111100100010110100000;
filter5[10][983] = 35'b11111100001110001000001011000100000;
filter5[10][984] = 35'b00000000100010000101000001001111000;
filter5[10][985] = 35'b11111111111110010101001000011010010;
filter5[10][986] = 35'b00000000011011011100000101111001100;
filter5[10][987] = 35'b11111101011000110001101100100100000;
filter5[10][988] = 35'b11111111010110110101011101111011000;
filter5[10][989] = 35'b11111101111111110111110000111100000;
filter5[10][990] = 35'b11111110110001111010110101110110000;
filter5[10][991] = 35'b11111111111001010000101010000111001;
filter5[10][992] = 35'b00000111010010010110001000111000000;
filter5[10][993] = 35'b11111110101001101100000010110000000;
filter5[10][994] = 35'b00000010110111011111111010000100000;
filter5[10][995] = 35'b11111110010100100101110110101100000;
filter5[10][996] = 35'b00000010000111010110100011100100000;
filter5[10][997] = 35'b00000010000011101001011001000000000;
filter5[10][998] = 35'b00000001010011100011101001000010000;
filter5[10][999] = 35'b11111100011010111110011001001000000;
filter5[10][1000] = 35'b11111010010100001011111101000000000;
filter5[10][1001] = 35'b11111110111111111110000001111000000;
filter5[10][1002] = 35'b11111110011001111001100001001010000;
filter5[10][1003] = 35'b11111010101101001011001001110000000;
filter5[10][1004] = 35'b11111011011101101011110111000000000;
filter5[10][1005] = 35'b11111101101111001101100001000100000;
filter5[10][1006] = 35'b00000110110001001100111011111000000;
filter5[10][1007] = 35'b00000110111100111000101000000000000;
filter5[10][1008] = 35'b00000010110111011111000011100100000;
filter5[10][1009] = 35'b11111111111010110010001001001100000;
filter5[10][1010] = 35'b11111000001110100101010110110000000;
filter5[10][1011] = 35'b11111111100101100101111001101000000;
filter5[10][1012] = 35'b11111101110011111010110000101000000;
filter5[10][1013] = 35'b11111101001110000110011110110000000;
filter5[10][1014] = 35'b00000101010010100010110001100000000;
filter5[10][1015] = 35'b00000000001010101000110011100011100;
filter5[10][1016] = 35'b00000000001101110111010010001110100;
filter5[10][1017] = 35'b00000100111011011111110000010000000;
filter5[10][1018] = 35'b11111010000110010111001000001000000;
filter5[10][1019] = 35'b00000111001010100001001111100000000;
filter5[10][1020] = 35'b00000110001011110100110110001000000;
filter5[10][1021] = 35'b00001111111100010000000011100000000;
filter5[10][1022] = 35'b00001100100100110010001000000000000;
filter5[10][1023] = 35'b00000111011011000101001111001000000;
bias5[0] = 35'b00000000100111110010101100010001000;
bias5[1] = 35'b11111111110001101011001010010100010;
bias5[2] = 35'b00000001011100100001010010000100000;
bias5[3] = 35'b11111001010010111111010001011000000;
bias5[4] = 35'b11111011000010010011011001010000000;
bias5[5] = 35'b11111100111010100101110000011000000;
bias5[6] = 35'b11111100000111110011010111100100000;
bias5[7] = 35'b11111110010000101001110011111000000;
bias5[8] = 35'b11111100100111011000011100010000000;
bias5[9] = 35'b11111000011001010101110101101000000;
bias5[10] = 35'b00000110000010011110011011010000000;

//==============================================================

//vmem_in[0][0][0]=0;
////        for(i=0;i<4;i++)
////        for(j=0;j<64;j++)
////        for(k=0;k<64;k++)
////        vmem_in[i][j][k]=0;
        
//         for(i=0;i<8;i++)
//        for(j=0;j<32;j++)
//        for(k=0;k<32;k++)
//        vmem_in2[i][j][k]=0;
        
//        for(i=0;i<8;i++)
//        for(j=0;j<16;j++)
//        for(k=0;k<16;k++) 
//        vmem_in3[i][j][k]=0;
        
//        for(i=0;i<16;i++)
//        for(j=0;j<8;j++)
//        for(k=0;k<8;k++) 
//        vmem_in4[i][j][k]=0;
        

  
        for (t=1;t<=3;t++) begin
       go=1;
       #120 $display("gotcha %0t",$time);
       
        if(t>1) begin
//        $display("yes, here %d",t);
        for(i=0;i<11;i++) begin 
        pred_in[i]=pred_out[i];
        $display("%d", pred_in[i]);
        end
        
         for(i=0;i<4;i++)
        for(j=0;j<64;j++)
        for(k=0;k<64;k++)
        vmem_in[i][j][k]=vmem_out[i][j][k];
        
         for(i=0;i<8;i++)
        for(j=0;j<32;j++)
        for(k=0;k<32;k++)
        vmem_in2[i][j][k]=vmem_out2[i][j][k];
        
        for(i=0;i<8;i++)
        for(j=0;j<16;j++)
        for(k=0;k<16;k++) 
        vmem_in3[i][j][k]=vmem_out3[i][j][k];
        
        for(i=0;i<16;i++)
        for(j=0;j<8;j++)
        for(k=0;k<8;k++) 
        vmem_in4[i][j][k]=vmem_out4[i][j][k];
        
        for(i=0;i<11;i++)
        vmem_in5[i]=vmem_out5[i];
           end
           
        else begin
        $display("t %d",t);
        for(i=0;i<11;i++) begin
        pred_in[i]=0;
        $display("pred in %d",pred_in[i]);
        end
        
         for(i=0;i<4;i++)
        for(j=0;j<64;j++)
        for(k=0;k<64;k++)
        vmem_in[i][j][k]=34'b0;
        
         for(i=0;i<8;i++)
        for(j=0;j<32;j++)
        for(k=0;k<32;k++)
        vmem_in2[i][j][k]=34'b0;
        
        for(i=0;i<8;i++)
        for(j=0;j<16;j++)
        for(k=0;k<16;k++) 
        vmem_in3[i][j][k]=34'b0;
        
        for(i=0;i<16;i++)
        for(j=0;j<8;j++)
        for(k=0;k<8;k++) 
        vmem_in4[i][j][k]=34'b0;
        
        for(i=0;i<11;i++)
        vmem_in5[i]=34'b0;
           end
//        #80 $display("gotcha %0t",$time); 

//    $display("pred_out %d",pred_out[0]);
        for (int w=0;w<2;w++) begin 
        for(int i = 0; i < 128; i++) begin
        for(int j = 0; j < 128; j++) begin
//        if(!$feof(fd)) begin
//////        in[w][i][j] = $fread(weight,fd);
//            $fscanf(fd,"%b",reg1);
//            in[w][i][j]=reg1[34:10];
//////            $display("input is %b",in[w][i][j]);
//       end
//       else
         in[w][i][j] = j-i;
//         $display("input is %b",in[w][i][j]);
//         in[1][i][j] = i;
//         $display ("vmemout %d %d",vmem_in[0][i][j],vmem_out[0][i][j]);
        end
        end
        end
//       #80 $display("gotcha");                 
        end
        
//        if (t>=3)
//        for(int i=0;i<11;i++)
//        $display("%d",pred_out[i]);
    end
    

    initial begin
//    go=0;
#120 clock=0;
forever #10 clock=~clock;
end

    
    initial begin
    reset=1;
    #3 reset=0;
//    for (int i=0;i<=2;i+=1) begin
//        for (int j=0;j<=2;j+=1) begin
//            #2 filter[i][j]=j;
//            end
//            end
        
//     for (int i=0;i<=7;i+=1)
//        for (int j=0;j<=7;j+=1) begin
//            in[i][j]=j;
//$display ("tbtb filter is %d",in[i][j]);
//        end

    #500 $finish;
    end
//    convo c1(clock,reset,bias,in,filter,out);

//generate 
//genvar i,j,k;
//for (i=0;i<150;i++)
layer1 l1(go,clock,reset,bias,bias2,bias3,bias4,bias5,in,filter,filter2,filter3,filter4,filter5,vmem_in,vmem_in2,vmem_in3,vmem_in4,vmem_in5, pred_in, vmem_out,vmem_out2,vmem_out3,vmem_out4,vmem_out5, pred_out);
//endgenerate
endmodule
